module CounterHsk(
  input   clock,
  input   reset,
  input   io_validPre,
  output  io_readyPre,
  output  io_validNxt,
  input   io_readyNxt,
  input   io_lastPre,
  output  io_lastNxt,
  output  io_regen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] counter; // @[Reg.scala 28:20]
  wire  _counterEn_T = io_validNxt & io_readyNxt; // @[counterhsk.scala 30:29]
  wire  counterEn = io_validNxt & io_readyNxt | io_regen; // @[counterhsk.scala 30:41]
  wire  _counterNxt_T = counter == 3'h4; // @[counterhsk.scala 25:16]
  wire  _counterNxt_T_1 = io_validPre & io_readyPre; // @[counterhsk.scala 26:24]
  wire [2:0] _counterNxt_T_4 = counter + 3'h1; // @[counterhsk.scala 27:16]
  wire  _io_regen_T_1 = counter == 3'h0; // @[counterhsk.scala 29:53]
  wire  _io_lastNxt_T_1 = io_validPre & io_validNxt & io_regen; // @[counterhsk.scala 33:69]
  reg  io_lastNxt_r; // @[Reg.scala 28:20]
  assign io_readyPre = _io_regen_T_1 | _counterEn_T; // @[counterhsk.scala 31:52]
  assign io_validNxt = counter == 3'h4; // @[counterhsk.scala 32:28]
  assign io_lastNxt = io_lastNxt_r; // @[counterhsk.scala 33:16]
  assign io_regen = _counterNxt_T_1 | ~(counter == 3'h0 | _counterNxt_T); // @[counterhsk.scala 29:41]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      counter <= 3'h0; // @[counterhsk.scala 24:22 26:12]
    end else if (counterEn) begin // @[Reg.scala 28:20]
      if (_counterNxt_T) begin
        if (io_validPre & io_readyPre) begin
          counter <= 3'h1;
        end else begin
          counter <= 3'h0;
        end
      end else begin
        counter <= _counterNxt_T_4;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      io_lastNxt_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (_io_lastNxt_T_1) begin // @[Reg.scala 28:20]
      io_lastNxt_r <= io_lastPre;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  io_lastNxt_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    counter = 3'h0;
  end
  if (reset) begin
    io_lastNxt_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Multiply(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [7:0]  io_input_bits_x_0,
  input  [7:0]  io_input_bits_x_1,
  input         io_input_bits_last,
  input         io_output_ready,
  output        io_output_valid,
  output [19:0] io_output_bits_x_0,
  output        io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  counterHsk_clock; // @[multiply.scala 20:28]
  wire  counterHsk_reset; // @[multiply.scala 20:28]
  wire  counterHsk_io_validPre; // @[multiply.scala 20:28]
  wire  counterHsk_io_readyPre; // @[multiply.scala 20:28]
  wire  counterHsk_io_validNxt; // @[multiply.scala 20:28]
  wire  counterHsk_io_readyNxt; // @[multiply.scala 20:28]
  wire  counterHsk_io_lastPre; // @[multiply.scala 20:28]
  wire  counterHsk_io_lastNxt; // @[multiply.scala 20:28]
  wire  counterHsk_io_regen; // @[multiply.scala 20:28]
  reg [7:0] in0; // @[Reg.scala 16:16]
  wire  _in0Nxt_T = io_input_valid & io_input_ready; // @[multiply.scala 31:33]
  wire [9:0] _in0Nxt_T_1 = {$signed(io_input_bits_x_0), 2'h0}; // @[multiply.scala 31:68]
  wire [9:0] _in0Nxt_T_2 = {$signed(in0), 2'h0}; // @[multiply.scala 31:76]
  wire [9:0] _in0Nxt_T_3 = io_input_valid & io_input_ready ? $signed(_in0Nxt_T_1) : $signed(_in0Nxt_T_2); // @[multiply.scala 31:18]
  wire [7:0] in0Nxt = _in0Nxt_T_3[7:0]; // @[multiply.scala 28:22 31:12]
  wire  _in1_T_1 = _in0Nxt_T & counterHsk_io_regen; // @[multiply.scala 30:74]
  reg [7:0] in1; // @[Reg.scala 16:16]
  wire [7:0] in1Inc = _in0Nxt_T ? $signed(io_input_bits_x_1) : $signed(in1); // @[multiply.scala 32:21]
  reg [15:0] out0; // @[Reg.scala 16:16]
  wire [2:0] out0IncMux = _in0Nxt_T ? io_input_bits_x_0[7:5] : in0[7:5]; // @[multiply.scala 38:25]
  wire [7:0] _out0Inc_T_13 = 8'sh0 - $signed(in1Inc); // @[multiply.scala 42:38]
  wire [8:0] _GEN_4 = {{1{in1Inc[7]}},in1Inc}; // @[multiply.scala 43:62]
  wire [8:0] _out0Inc_T_20 = 9'sh0 - $signed(_GEN_4); // @[multiply.scala 43:62]
  wire [8:0] _out0Inc_T_21 = out0IncMux == 3'h5 | out0IncMux == 3'h6 ? $signed(_out0Inc_T_20) : $signed(9'sh0); // @[multiply.scala 43:12]
  wire [8:0] _out0Inc_T_22 = out0IncMux == 3'h4 ? $signed({$signed(_out0Inc_T_13), 1'h0}) : $signed(_out0Inc_T_21); // @[multiply.scala 42:12]
  wire [8:0] _out0Inc_T_23 = out0IncMux == 3'h3 ? $signed({$signed(in1Inc), 1'h0}) : $signed(_out0Inc_T_22); // @[multiply.scala 41:12]
  wire [8:0] _out0Inc_T_24 = out0IncMux == 3'h1 | out0IncMux == 3'h2 ? $signed({{1{in1Inc[7]}},in1Inc}) : $signed(
    _out0Inc_T_23); // @[multiply.scala 40:12]
  wire [8:0] _out0Inc_T_25 = out0IncMux == 3'h0 | out0IncMux == 3'h7 ? $signed(9'sh0) : $signed(_out0Inc_T_24); // @[multiply.scala 39:19]
  wire [15:0] out0Inc = {{7{_out0Inc_T_25[8]}},_out0Inc_T_25}; // @[multiply.scala 35:23 39:13]
  wire [17:0] _GEN_5 = {$signed(out0), 2'h0}; // @[multiply.scala 37:92]
  wire [17:0] _GEN_6 = {{2{out0Inc[15]}},out0Inc}; // @[multiply.scala 37:92]
  wire [17:0] _out0Nxt_T_4 = $signed(_GEN_5) + $signed(_GEN_6); // @[multiply.scala 37:92]
  wire [17:0] _out0Nxt_T_5 = _in0Nxt_T ? $signed({{2{out0Inc[15]}},out0Inc}) : $signed(_out0Nxt_T_4); // @[multiply.scala 37:19]
  wire [15:0] out0Nxt = _out0Nxt_T_5[15:0]; // @[multiply.scala 34:23 37:13]
  CounterHsk counterHsk ( // @[multiply.scala 20:28]
    .clock(counterHsk_clock),
    .reset(counterHsk_reset),
    .io_validPre(counterHsk_io_validPre),
    .io_readyPre(counterHsk_io_readyPre),
    .io_validNxt(counterHsk_io_validNxt),
    .io_readyNxt(counterHsk_io_readyNxt),
    .io_lastPre(counterHsk_io_lastPre),
    .io_lastNxt(counterHsk_io_lastNxt),
    .io_regen(counterHsk_io_regen)
  );
  assign io_input_ready = counterHsk_io_readyPre; // @[multiply.scala 22:20]
  assign io_output_valid = counterHsk_io_validNxt; // @[multiply.scala 23:21]
  assign io_output_bits_x_0 = {{4{out0[15]}},out0}; // @[multiply.scala 46:25]
  assign io_output_bits_last = counterHsk_io_lastNxt; // @[multiply.scala 26:25]
  assign counterHsk_clock = clock;
  assign counterHsk_reset = reset;
  assign counterHsk_io_validPre = io_input_valid; // @[multiply.scala 21:28]
  assign counterHsk_io_readyNxt = io_output_ready; // @[multiply.scala 24:28]
  assign counterHsk_io_lastPre = io_input_bits_last; // @[multiply.scala 25:27]
  always @(posedge clock) begin
    if (counterHsk_io_regen) begin // @[Reg.scala 17:18]
      in0 <= in0Nxt; // @[Reg.scala 17:22]
    end
    if (_in1_T_1) begin // @[Reg.scala 17:18]
      in1 <= io_input_bits_x_1; // @[Reg.scala 17:22]
    end
    if (counterHsk_io_regen) begin // @[Reg.scala 17:18]
      out0 <= out0Nxt; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  in1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  out0 = _RAND_2[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineHsk(
  input   clock,
  input   reset,
  input   io_validPre,
  output  io_readyPre,
  input   io_lastPre,
  output  io_validNxt,
  input   io_readyNxt,
  output  io_regen_0,
  output  io_lastNxt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  valid_1_r; // @[Reg.scala 28:20]
  wire  ready_0 = io_readyNxt | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  reg  last_1_r; // @[Reg.scala 28:20]
  assign io_readyPre = io_readyNxt | ~valid_1_r; // @[pipelinehsk.scala 24:32]
  assign io_validNxt = valid_1_r; // @[pipelinehsk.scala 17:21 22:20]
  assign io_regen_0 = io_validPre & ready_0; // @[pipelinehsk.scala 25:33]
  assign io_lastNxt = last_1_r; // @[pipelinehsk.scala 19:20 23:19]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      valid_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (ready_0) begin // @[Reg.scala 28:20]
      valid_1_r <= io_validPre;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      last_1_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_regen_0) begin // @[Reg.scala 28:20]
      last_1_r <= io_lastPre;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_1_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  last_1_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid_1_r = 1'h0;
  end
  if (reset) begin
    last_1_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Adder2to1(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [19:0] io_input_bits_x_0,
  input  [19:0] io_input_bits_x_1,
  input         io_input_bits_last,
  input         io_output_ready,
  output        io_output_valid,
  output [19:0] io_output_bits_x_0,
  output        io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  hsk_clock; // @[adder2to1.scala 26:25]
  wire  hsk_reset; // @[adder2to1.scala 26:25]
  wire  hsk_io_validPre; // @[adder2to1.scala 26:25]
  wire  hsk_io_readyPre; // @[adder2to1.scala 26:25]
  wire  hsk_io_lastPre; // @[adder2to1.scala 26:25]
  wire  hsk_io_validNxt; // @[adder2to1.scala 26:25]
  wire  hsk_io_readyNxt; // @[adder2to1.scala 26:25]
  wire  hsk_io_regen_0; // @[adder2to1.scala 26:25]
  wire  hsk_io_lastNxt; // @[adder2to1.scala 26:25]
  wire [19:0] sum_0 = $signed(io_input_bits_x_0) + $signed(io_input_bits_x_1); // @[adder2to1.scala 23:69]
  reg [19:0] r_0; // @[Reg.scala 16:16]
  PipelineHsk hsk ( // @[adder2to1.scala 26:25]
    .clock(hsk_clock),
    .reset(hsk_reset),
    .io_validPre(hsk_io_validPre),
    .io_readyPre(hsk_io_readyPre),
    .io_lastPre(hsk_io_lastPre),
    .io_validNxt(hsk_io_validNxt),
    .io_readyNxt(hsk_io_readyNxt),
    .io_regen_0(hsk_io_regen_0),
    .io_lastNxt(hsk_io_lastNxt)
  );
  assign io_input_ready = hsk_io_readyPre; // @[adder2to1.scala 28:24]
  assign io_output_valid = hsk_io_validNxt; // @[adder2to1.scala 29:25]
  assign io_output_bits_x_0 = r_0; // @[adder2to1.scala 33:26]
  assign io_output_bits_last = hsk_io_lastNxt; // @[adder2to1.scala 32:29]
  assign hsk_clock = clock;
  assign hsk_reset = reset;
  assign hsk_io_validPre = io_input_valid; // @[adder2to1.scala 27:25]
  assign hsk_io_lastPre = io_input_bits_last; // @[adder2to1.scala 31:24]
  assign hsk_io_readyNxt = io_output_ready; // @[adder2to1.scala 30:25]
  always @(posedge clock) begin
    if (hsk_io_regen_0) begin // @[Reg.scala 17:18]
      r_0 <= sum_0; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_0 = _RAND_0[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Hsknto1(
  output        io_input_0_ready,
  input         io_input_0_valid,
  input  [19:0] io_input_0_bits_x_0,
  output        io_input_1_ready,
  input         io_input_1_valid,
  input  [19:0] io_input_1_bits_x_0,
  input         io_input_1_bits_last,
  input         io_output_ready,
  output        io_output_valid,
  output [19:0] io_output_bits_0_x_0,
  output [19:0] io_output_bits_1_x_0,
  output        io_output_bits_1_last
);
  assign io_input_0_ready = io_output_ready & (~io_input_0_valid | io_input_1_valid); // @[hsknto1.scala 14:73]
  assign io_input_1_ready = io_output_ready & (~io_input_1_valid | io_input_0_valid); // @[hsknto1.scala 14:73]
  assign io_output_valid = io_input_0_valid & io_input_1_valid; // @[hsknto1.scala 12:58]
  assign io_output_bits_0_x_0 = io_input_0_bits_x_0; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_0 = io_input_1_bits_x_0; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_last = io_input_1_bits_last; // @[hsknto1.scala 13:55]
endmodule
module Accumulator2to1(
  input         clock,
  input         reset,
  output        io_input_ready,
  input         io_input_valid,
  input  [19:0] io_input_bits_x_0,
  input         io_input_bits_last,
  output        io_output_valid,
  output [19:0] io_output_bits_x_0,
  output        io_output_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _io_output_bits_last_T = io_input_valid & io_input_ready; // @[accumulator2to1.scala 17:77]
  reg  io_output_bits_last_r; // @[Reg.scala 28:20]
  reg [19:0] io_output_bits_x_0_r; // @[Reg.scala 28:20]
  wire [19:0] _sumNxt_T_2 = $signed(io_output_bits_x_0) + $signed(io_input_bits_x_0); // @[accumulator2to1.scala 19:79]
  assign io_input_ready = 1'h1; // @[accumulator2to1.scala 15:20]
  assign io_output_valid = io_output_bits_last; // @[accumulator2to1.scala 20:21]
  assign io_output_bits_x_0 = io_output_bits_x_0_r; // @[accumulator2to1.scala 18:25]
  assign io_output_bits_last = io_output_bits_last_r; // @[accumulator2to1.scala 17:25]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      io_output_bits_last_r <= 1'h0; // @[Reg.scala 29:22]
    end else if (_io_output_bits_last_T) begin // @[Reg.scala 28:20]
      io_output_bits_last_r <= io_input_bits_last;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      io_output_bits_x_0_r <= 20'sh0; // @[accumulator2to1.scala 19:18]
    end else if (_io_output_bits_last_T) begin // @[Reg.scala 28:20]
      if (io_output_bits_last) begin
        io_output_bits_x_0_r <= io_input_bits_x_0;
      end else begin
        io_output_bits_x_0_r <= _sumNxt_T_2;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_output_bits_last_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_output_bits_x_0_r = _RAND_1[19:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    io_output_bits_last_r = 1'h0;
  end
  if (reset) begin
    io_output_bits_x_0_r = 20'sh0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Arbiter1ton(
  output        io_input_ready,
  input         io_input_valid,
  input  [19:0] io_input_bits_x_0,
  input         io_input_bits_last,
  input         io_sel,
  input         io_output_0_ready,
  output        io_output_0_valid,
  output [19:0] io_output_0_bits_x_0,
  output        io_output_0_bits_last,
  output        io_output_1_valid,
  output [19:0] io_output_1_bits_x_0,
  output        io_output_1_bits_last
);
  assign io_input_ready = io_sel | io_output_0_ready; // @[arbiter1ton.scala 16:{20,20}]
  assign io_output_0_valid = ~io_sel & io_input_valid; // @[arbiter1ton.scala 18:44]
  assign io_output_0_bits_x_0 = io_input_bits_x_0; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_last = io_input_bits_last; // @[arbiter1ton.scala 19:26]
  assign io_output_1_valid = io_sel & io_input_valid; // @[arbiter1ton.scala 18:44]
  assign io_output_1_bits_x_0 = io_input_bits_x_0; // @[arbiter1ton.scala 19:26]
  assign io_output_1_bits_last = io_input_bits_last; // @[arbiter1ton.scala 19:26]
endmodule
module Arbiternto1(
  output        io_input_0_ready,
  input         io_input_0_valid,
  input  [19:0] io_input_0_bits_x_0,
  input         io_input_0_bits_last,
  input         io_input_1_valid,
  input  [19:0] io_input_1_bits_x_0,
  input         io_input_1_bits_last,
  input         io_sel,
  input         io_output_ready,
  output        io_output_valid,
  output [19:0] io_output_bits_x_0,
  output        io_output_bits_last
);
  assign io_input_0_ready = ~io_sel & io_output_ready; // @[arbiternto1.scala 17:44]
  assign io_output_valid = io_sel ? io_input_1_valid : io_input_0_valid; // @[arbiternto1.scala 15:{21,21}]
  assign io_output_bits_x_0 = io_sel ? $signed(io_input_1_bits_x_0) : $signed(io_input_0_bits_x_0); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_last = io_sel ? io_input_1_bits_last : io_input_0_bits_last; // @[arbiternto1.scala 14:{20,20}]
endmodule
module Hsknto1_1(
  output       io_input_0_ready,
  input        io_input_0_valid,
  input  [7:0] io_input_0_bits_x_0,
  input        io_input_0_bits_last,
  output       io_input_1_ready,
  input        io_input_1_valid,
  input  [7:0] io_input_1_bits_x_0,
  input        io_input_1_bits_last,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_0_x_0,
  output       io_output_bits_0_last,
  output [7:0] io_output_bits_1_x_0,
  output       io_output_bits_1_last
);
  assign io_input_0_ready = io_output_ready & (~io_input_0_valid | io_input_1_valid); // @[hsknto1.scala 14:73]
  assign io_input_1_ready = io_output_ready & (~io_input_1_valid | io_input_0_valid); // @[hsknto1.scala 14:73]
  assign io_output_valid = io_input_0_valid & io_input_1_valid; // @[hsknto1.scala 12:58]
  assign io_output_bits_0_x_0 = io_input_0_bits_x_0; // @[hsknto1.scala 13:55]
  assign io_output_bits_0_last = io_input_0_bits_last; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_x_0 = io_input_1_bits_x_0; // @[hsknto1.scala 13:55]
  assign io_output_bits_1_last = io_input_1_bits_last; // @[hsknto1.scala 13:55]
endmodule
module Hsk1ton(
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_0_x_0,
  input  [7:0] io_input_bits_0_x_1,
  input        io_input_bits_0_last,
  input  [7:0] io_input_bits_1_x_0,
  input  [7:0] io_input_bits_1_x_1,
  input        io_input_bits_1_last,
  input  [7:0] io_input_bits_2_x_0,
  input  [7:0] io_input_bits_2_x_1,
  input        io_input_bits_2_last,
  input        io_output_0_ready,
  output       io_output_0_valid,
  output [7:0] io_output_0_bits_x_0,
  output [7:0] io_output_0_bits_x_1,
  output       io_output_0_bits_last,
  input        io_output_1_ready,
  output       io_output_1_valid,
  output [7:0] io_output_1_bits_x_0,
  output [7:0] io_output_1_bits_x_1,
  output       io_output_1_bits_last,
  input        io_output_2_ready,
  output       io_output_2_valid,
  output [7:0] io_output_2_bits_x_0,
  output [7:0] io_output_2_bits_x_1,
  output       io_output_2_bits_last
);
  wire  _io_input_ready_T_1 = io_output_0_ready & io_output_1_ready; // @[hsk1ton.scala 12:58]
  wire  _io_output_0_valid_T_6 = io_output_1_ready & io_output_2_ready; // @[hsk1ton.scala 15:72]
  wire  _io_output_1_valid_T_6 = io_output_0_ready & io_output_2_ready; // @[hsk1ton.scala 15:72]
  assign io_input_ready = io_output_0_ready & io_output_1_ready & io_output_2_ready; // @[hsk1ton.scala 12:58]
  assign io_output_0_valid = io_input_valid & (~io_output_0_ready | _io_output_0_valid_T_6); // @[hsk1ton.scala 14:72]
  assign io_output_0_bits_x_0 = io_input_bits_0_x_0; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_x_1 = io_input_bits_0_x_1; // @[hsk1ton.scala 13:54]
  assign io_output_0_bits_last = io_input_bits_0_last; // @[hsk1ton.scala 13:54]
  assign io_output_1_valid = io_input_valid & (~io_output_1_ready | _io_output_1_valid_T_6); // @[hsk1ton.scala 14:72]
  assign io_output_1_bits_x_0 = io_input_bits_1_x_0; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_x_1 = io_input_bits_1_x_1; // @[hsk1ton.scala 13:54]
  assign io_output_1_bits_last = io_input_bits_1_last; // @[hsk1ton.scala 13:54]
  assign io_output_2_valid = io_input_valid & (~io_output_2_ready | _io_input_ready_T_1); // @[hsk1ton.scala 14:72]
  assign io_output_2_bits_x_0 = io_input_bits_2_x_0; // @[hsk1ton.scala 13:54]
  assign io_output_2_bits_x_1 = io_input_bits_2_x_1; // @[hsk1ton.scala 13:54]
  assign io_output_2_bits_last = io_input_bits_2_last; // @[hsk1ton.scala 13:54]
endmodule
module Arbiternto1_1(
  output       io_input_0_ready,
  input        io_input_0_valid,
  input  [7:0] io_input_0_bits_x_0,
  input        io_input_0_bits_last,
  input        io_sel,
  input        io_output_ready,
  output       io_output_valid,
  output [7:0] io_output_bits_x_0,
  output       io_output_bits_last
);
  assign io_input_0_ready = ~io_sel & io_output_ready; // @[arbiternto1.scala 17:44]
  assign io_output_valid = io_sel | io_input_0_valid; // @[arbiternto1.scala 15:{21,21}]
  assign io_output_bits_x_0 = io_sel ? $signed(8'sh0) : $signed(io_input_0_bits_x_0); // @[arbiternto1.scala 14:{20,20}]
  assign io_output_bits_last = io_sel ? 1'h0 : io_input_0_bits_last; // @[arbiternto1.scala 14:{20,20}]
endmodule
module Arbiter1ton_1(
  output       io_input_ready,
  input        io_input_valid,
  input  [7:0] io_input_bits_x_0,
  input  [7:0] io_input_bits_x_1,
  input        io_input_bits_last,
  input        io_sel,
  input        io_output_0_ready,
  output       io_output_0_valid,
  output [7:0] io_output_0_bits_x_0,
  output [7:0] io_output_0_bits_x_1,
  output       io_output_0_bits_last
);
  assign io_input_ready = io_sel | io_output_0_ready; // @[arbiter1ton.scala 16:{20,20}]
  assign io_output_0_valid = ~io_sel & io_input_valid; // @[arbiter1ton.scala 18:44]
  assign io_output_0_bits_x_0 = io_input_bits_x_0; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_x_1 = io_input_bits_x_1; // @[arbiter1ton.scala 19:26]
  assign io_output_0_bits_last = io_input_bits_last; // @[arbiter1ton.scala 19:26]
endmodule
module PECross(
  input         clock,
  input         reset,
  output        multiply_io_input_io_sumIn_ready,
  input         multiply_io_input_io_sumIn_valid,
  input  [19:0] multiply_io_input_io_sumIn_bits_x_0,
  input         multiply_io_input_io_sumIn_bits_last,
  input         multiply_io_input_io_sumOut_ready,
  output        multiply_io_input_io_sumOut_valid,
  output [19:0] multiply_io_input_io_sumOut_bits_x_0,
  output        multiply_io_input_io_sumOut_bits_last,
  input  [1:0]  multiply_io_input_io_statSel,
  input         multiply_io_input_io_weiEn,
  input         multiply_io_input_io_actEn,
  output        multiply_io_input_io_actIn_ready,
  input         multiply_io_input_io_actIn_valid,
  input  [7:0]  multiply_io_input_io_actIn_bits_x_0,
  input         multiply_io_input_io_actIn_bits_last,
  output        multiply_io_input_io_weiIn_ready,
  input         multiply_io_input_io_weiIn_valid,
  input  [7:0]  multiply_io_input_io_weiIn_bits_x_0,
  input         multiply_io_input_io_weiIn_bits_last,
  input         multiply_io_input_io_actOut_ready,
  output        multiply_io_input_io_actOut_valid,
  output [7:0]  multiply_io_input_io_actOut_bits_x_0,
  output        multiply_io_input_io_actOut_bits_last,
  input         multiply_io_input_io_weiOut_ready,
  output        multiply_io_input_io_weiOut_valid,
  output [7:0]  multiply_io_input_io_weiOut_bits_x_0,
  output        multiply_io_input_io_weiOut_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  multiply_clock; // @[penlr.scala 14:26]
  wire  multiply_reset; // @[penlr.scala 14:26]
  wire  multiply_io_input_ready; // @[penlr.scala 14:26]
  wire  multiply_io_input_valid; // @[penlr.scala 14:26]
  wire [7:0] multiply_io_input_bits_x_0; // @[penlr.scala 14:26]
  wire [7:0] multiply_io_input_bits_x_1; // @[penlr.scala 14:26]
  wire  multiply_io_input_bits_last; // @[penlr.scala 14:26]
  wire  multiply_io_output_ready; // @[penlr.scala 14:26]
  wire  multiply_io_output_valid; // @[penlr.scala 14:26]
  wire [19:0] multiply_io_output_bits_x_0; // @[penlr.scala 14:26]
  wire  multiply_io_output_bits_last; // @[penlr.scala 14:26]
  wire  adder_clock; // @[penlr.scala 17:23]
  wire  adder_reset; // @[penlr.scala 17:23]
  wire  adder_io_input_ready; // @[penlr.scala 17:23]
  wire  adder_io_input_valid; // @[penlr.scala 17:23]
  wire [19:0] adder_io_input_bits_x_0; // @[penlr.scala 17:23]
  wire [19:0] adder_io_input_bits_x_1; // @[penlr.scala 17:23]
  wire  adder_io_input_bits_last; // @[penlr.scala 17:23]
  wire  adder_io_output_ready; // @[penlr.scala 17:23]
  wire  adder_io_output_valid; // @[penlr.scala 17:23]
  wire [19:0] adder_io_output_bits_x_0; // @[penlr.scala 17:23]
  wire  adder_io_output_bits_last; // @[penlr.scala 17:23]
  wire  adderInHsk_io_input_0_ready; // @[penlr.scala 18:28]
  wire  adderInHsk_io_input_0_valid; // @[penlr.scala 18:28]
  wire [19:0] adderInHsk_io_input_0_bits_x_0; // @[penlr.scala 18:28]
  wire  adderInHsk_io_input_1_ready; // @[penlr.scala 18:28]
  wire  adderInHsk_io_input_1_valid; // @[penlr.scala 18:28]
  wire [19:0] adderInHsk_io_input_1_bits_x_0; // @[penlr.scala 18:28]
  wire  adderInHsk_io_input_1_bits_last; // @[penlr.scala 18:28]
  wire  adderInHsk_io_output_ready; // @[penlr.scala 18:28]
  wire  adderInHsk_io_output_valid; // @[penlr.scala 18:28]
  wire [19:0] adderInHsk_io_output_bits_0_x_0; // @[penlr.scala 18:28]
  wire [19:0] adderInHsk_io_output_bits_1_x_0; // @[penlr.scala 18:28]
  wire  adderInHsk_io_output_bits_1_last; // @[penlr.scala 18:28]
  wire  accumulator_clock; // @[pe.scala 19:29]
  wire  accumulator_reset; // @[pe.scala 19:29]
  wire  accumulator_io_input_ready; // @[pe.scala 19:29]
  wire  accumulator_io_input_valid; // @[pe.scala 19:29]
  wire [19:0] accumulator_io_input_bits_x_0; // @[pe.scala 19:29]
  wire  accumulator_io_input_bits_last; // @[pe.scala 19:29]
  wire  accumulator_io_output_valid; // @[pe.scala 19:29]
  wire [19:0] accumulator_io_output_bits_x_0; // @[pe.scala 19:29]
  wire  accumulator_io_output_bits_last; // @[pe.scala 19:29]
  wire  multiplyOutMux_io_input_ready; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_input_valid; // @[pe.scala 20:32]
  wire [19:0] multiplyOutMux_io_input_bits_x_0; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_input_bits_last; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_sel; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_output_0_ready; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_output_0_valid; // @[pe.scala 20:32]
  wire [19:0] multiplyOutMux_io_output_0_bits_x_0; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_output_0_bits_last; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_output_1_valid; // @[pe.scala 20:32]
  wire [19:0] multiplyOutMux_io_output_1_bits_x_0; // @[pe.scala 20:32]
  wire  multiplyOutMux_io_output_1_bits_last; // @[pe.scala 20:32]
  wire  sumOutMux_io_input_0_ready; // @[pe.scala 21:27]
  wire  sumOutMux_io_input_0_valid; // @[pe.scala 21:27]
  wire [19:0] sumOutMux_io_input_0_bits_x_0; // @[pe.scala 21:27]
  wire  sumOutMux_io_input_0_bits_last; // @[pe.scala 21:27]
  wire  sumOutMux_io_input_1_valid; // @[pe.scala 21:27]
  wire [19:0] sumOutMux_io_input_1_bits_x_0; // @[pe.scala 21:27]
  wire  sumOutMux_io_input_1_bits_last; // @[pe.scala 21:27]
  wire  sumOutMux_io_sel; // @[pe.scala 21:27]
  wire  sumOutMux_io_output_ready; // @[pe.scala 21:27]
  wire  sumOutMux_io_output_valid; // @[pe.scala 21:27]
  wire [19:0] sumOutMux_io_output_bits_x_0; // @[pe.scala 21:27]
  wire  sumOutMux_io_output_bits_last; // @[pe.scala 21:27]
  wire  actWeiInHsk_io_input_0_ready; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_input_0_valid; // @[pecross.scala 14:29]
  wire [7:0] actWeiInHsk_io_input_0_bits_x_0; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_input_0_bits_last; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_input_1_ready; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_input_1_valid; // @[pecross.scala 14:29]
  wire [7:0] actWeiInHsk_io_input_1_bits_x_0; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_input_1_bits_last; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_output_ready; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_output_valid; // @[pecross.scala 14:29]
  wire [7:0] actWeiInHsk_io_output_bits_0_x_0; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_output_bits_0_last; // @[pecross.scala 14:29]
  wire [7:0] actWeiInHsk_io_output_bits_1_x_0; // @[pecross.scala 14:29]
  wire  actWeiInHsk_io_output_bits_1_last; // @[pecross.scala 14:29]
  wire  multiplyInHsk_io_input_ready; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_input_valid; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_input_bits_0_x_0; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_input_bits_0_x_1; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_input_bits_0_last; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_input_bits_1_x_0; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_input_bits_1_x_1; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_input_bits_1_last; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_input_bits_2_x_0; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_input_bits_2_x_1; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_input_bits_2_last; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_0_ready; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_0_valid; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_output_0_bits_x_0; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_output_0_bits_x_1; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_0_bits_last; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_1_ready; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_1_valid; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_output_1_bits_x_0; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_output_1_bits_x_1; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_1_bits_last; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_2_ready; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_2_valid; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_output_2_bits_x_0; // @[pecross.scala 15:31]
  wire [7:0] multiplyInHsk_io_output_2_bits_x_1; // @[pecross.scala 15:31]
  wire  multiplyInHsk_io_output_2_bits_last; // @[pecross.scala 15:31]
  wire  weiInMux_io_input_0_ready; // @[pecross.scala 16:26]
  wire  weiInMux_io_input_0_valid; // @[pecross.scala 16:26]
  wire [7:0] weiInMux_io_input_0_bits_x_0; // @[pecross.scala 16:26]
  wire  weiInMux_io_input_0_bits_last; // @[pecross.scala 16:26]
  wire  weiInMux_io_sel; // @[pecross.scala 16:26]
  wire  weiInMux_io_output_ready; // @[pecross.scala 16:26]
  wire  weiInMux_io_output_valid; // @[pecross.scala 16:26]
  wire [7:0] weiInMux_io_output_bits_x_0; // @[pecross.scala 16:26]
  wire  weiInMux_io_output_bits_last; // @[pecross.scala 16:26]
  wire  actInMux_io_input_0_ready; // @[pecross.scala 17:26]
  wire  actInMux_io_input_0_valid; // @[pecross.scala 17:26]
  wire [7:0] actInMux_io_input_0_bits_x_0; // @[pecross.scala 17:26]
  wire  actInMux_io_input_0_bits_last; // @[pecross.scala 17:26]
  wire  actInMux_io_sel; // @[pecross.scala 17:26]
  wire  actInMux_io_output_ready; // @[pecross.scala 17:26]
  wire  actInMux_io_output_valid; // @[pecross.scala 17:26]
  wire [7:0] actInMux_io_output_bits_x_0; // @[pecross.scala 17:26]
  wire  actInMux_io_output_bits_last; // @[pecross.scala 17:26]
  wire  multiplyInMux_io_input_ready; // @[pecross.scala 18:31]
  wire  multiplyInMux_io_input_valid; // @[pecross.scala 18:31]
  wire [7:0] multiplyInMux_io_input_bits_x_0; // @[pecross.scala 18:31]
  wire [7:0] multiplyInMux_io_input_bits_x_1; // @[pecross.scala 18:31]
  wire  multiplyInMux_io_input_bits_last; // @[pecross.scala 18:31]
  wire  multiplyInMux_io_sel; // @[pecross.scala 18:31]
  wire  multiplyInMux_io_output_0_ready; // @[pecross.scala 18:31]
  wire  multiplyInMux_io_output_0_valid; // @[pecross.scala 18:31]
  wire [7:0] multiplyInMux_io_output_0_bits_x_0; // @[pecross.scala 18:31]
  wire [7:0] multiplyInMux_io_output_0_bits_x_1; // @[pecross.scala 18:31]
  wire  multiplyInMux_io_output_0_bits_last; // @[pecross.scala 18:31]
  wire  actOutMux_io_input_ready; // @[pecross.scala 19:27]
  wire  actOutMux_io_input_valid; // @[pecross.scala 19:27]
  wire [7:0] actOutMux_io_input_bits_x_0; // @[pecross.scala 19:27]
  wire [7:0] actOutMux_io_input_bits_x_1; // @[pecross.scala 19:27]
  wire  actOutMux_io_input_bits_last; // @[pecross.scala 19:27]
  wire  actOutMux_io_sel; // @[pecross.scala 19:27]
  wire  actOutMux_io_output_0_ready; // @[pecross.scala 19:27]
  wire  actOutMux_io_output_0_valid; // @[pecross.scala 19:27]
  wire [7:0] actOutMux_io_output_0_bits_x_0; // @[pecross.scala 19:27]
  wire [7:0] actOutMux_io_output_0_bits_x_1; // @[pecross.scala 19:27]
  wire  actOutMux_io_output_0_bits_last; // @[pecross.scala 19:27]
  wire  weiOutMux_io_input_ready; // @[pecross.scala 20:27]
  wire  weiOutMux_io_input_valid; // @[pecross.scala 20:27]
  wire [7:0] weiOutMux_io_input_bits_x_0; // @[pecross.scala 20:27]
  wire [7:0] weiOutMux_io_input_bits_x_1; // @[pecross.scala 20:27]
  wire  weiOutMux_io_input_bits_last; // @[pecross.scala 20:27]
  wire  weiOutMux_io_sel; // @[pecross.scala 20:27]
  wire  weiOutMux_io_output_0_ready; // @[pecross.scala 20:27]
  wire  weiOutMux_io_output_0_valid; // @[pecross.scala 20:27]
  wire [7:0] weiOutMux_io_output_0_bits_x_0; // @[pecross.scala 20:27]
  wire [7:0] weiOutMux_io_output_0_bits_x_1; // @[pecross.scala 20:27]
  wire  weiOutMux_io_output_0_bits_last; // @[pecross.scala 20:27]
  wire  adderInMux_io_input_0_ready; // @[pecross.scala 21:28]
  wire  adderInMux_io_input_0_valid; // @[pecross.scala 21:28]
  wire [19:0] adderInMux_io_input_0_bits_x_0; // @[pecross.scala 21:28]
  wire  adderInMux_io_input_0_bits_last; // @[pecross.scala 21:28]
  wire  adderInMux_io_input_1_valid; // @[pecross.scala 21:28]
  wire [19:0] adderInMux_io_input_1_bits_x_0; // @[pecross.scala 21:28]
  wire  adderInMux_io_input_1_bits_last; // @[pecross.scala 21:28]
  wire  adderInMux_io_sel; // @[pecross.scala 21:28]
  wire  adderInMux_io_output_ready; // @[pecross.scala 21:28]
  wire  adderInMux_io_output_valid; // @[pecross.scala 21:28]
  wire [19:0] adderInMux_io_output_bits_x_0; // @[pecross.scala 21:28]
  wire  adderInMux_io_output_bits_last; // @[pecross.scala 21:28]
  wire  actOutHsk_clock; // @[pecross.scala 47:27]
  wire  actOutHsk_reset; // @[pecross.scala 47:27]
  wire  actOutHsk_io_validPre; // @[pecross.scala 47:27]
  wire  actOutHsk_io_readyPre; // @[pecross.scala 47:27]
  wire  actOutHsk_io_lastPre; // @[pecross.scala 47:27]
  wire  actOutHsk_io_validNxt; // @[pecross.scala 47:27]
  wire  actOutHsk_io_readyNxt; // @[pecross.scala 47:27]
  wire  actOutHsk_io_regen_0; // @[pecross.scala 47:27]
  wire  actOutHsk_io_lastNxt; // @[pecross.scala 47:27]
  wire  weiOutHsk_clock; // @[pecross.scala 58:27]
  wire  weiOutHsk_reset; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_validPre; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_readyPre; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_lastPre; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_validNxt; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_readyNxt; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_regen_0; // @[pecross.scala 58:27]
  wire  weiOutHsk_io_lastNxt; // @[pecross.scala 58:27]
  wire  _weiOut_T = multiply_io_input_io_statSel == 2'h1; // @[pe.scala 15:62]
  wire  _weiOut_T_1 = multiply_io_input_io_statSel == 2'h1 & multiply_io_input_io_weiEn; // @[pe.scala 15:74]
  wire  _multiplyOutMux_io_sel_T = multiply_io_input_io_statSel == 2'h2; // @[pe.scala 22:41]
  reg [7:0] io_actOut_bits_x_0_r; // @[Reg.scala 16:16]
  reg [7:0] io_weiOut_bits_x_0_r; // @[Reg.scala 16:16]
  wire  _actInMux_io_sel_T_1 = ~multiply_io_input_io_weiEn; // @[pecross.scala 68:49]
  Multiply multiply ( // @[penlr.scala 14:26]
    .clock(multiply_clock),
    .reset(multiply_reset),
    .io_input_ready(multiply_io_input_ready),
    .io_input_valid(multiply_io_input_valid),
    .io_input_bits_x_0(multiply_io_input_bits_x_0),
    .io_input_bits_x_1(multiply_io_input_bits_x_1),
    .io_input_bits_last(multiply_io_input_bits_last),
    .io_output_ready(multiply_io_output_ready),
    .io_output_valid(multiply_io_output_valid),
    .io_output_bits_x_0(multiply_io_output_bits_x_0),
    .io_output_bits_last(multiply_io_output_bits_last)
  );
  Adder2to1 adder ( // @[penlr.scala 17:23]
    .clock(adder_clock),
    .reset(adder_reset),
    .io_input_ready(adder_io_input_ready),
    .io_input_valid(adder_io_input_valid),
    .io_input_bits_x_0(adder_io_input_bits_x_0),
    .io_input_bits_x_1(adder_io_input_bits_x_1),
    .io_input_bits_last(adder_io_input_bits_last),
    .io_output_ready(adder_io_output_ready),
    .io_output_valid(adder_io_output_valid),
    .io_output_bits_x_0(adder_io_output_bits_x_0),
    .io_output_bits_last(adder_io_output_bits_last)
  );
  Hsknto1 adderInHsk ( // @[penlr.scala 18:28]
    .io_input_0_ready(adderInHsk_io_input_0_ready),
    .io_input_0_valid(adderInHsk_io_input_0_valid),
    .io_input_0_bits_x_0(adderInHsk_io_input_0_bits_x_0),
    .io_input_1_ready(adderInHsk_io_input_1_ready),
    .io_input_1_valid(adderInHsk_io_input_1_valid),
    .io_input_1_bits_x_0(adderInHsk_io_input_1_bits_x_0),
    .io_input_1_bits_last(adderInHsk_io_input_1_bits_last),
    .io_output_ready(adderInHsk_io_output_ready),
    .io_output_valid(adderInHsk_io_output_valid),
    .io_output_bits_0_x_0(adderInHsk_io_output_bits_0_x_0),
    .io_output_bits_1_x_0(adderInHsk_io_output_bits_1_x_0),
    .io_output_bits_1_last(adderInHsk_io_output_bits_1_last)
  );
  Accumulator2to1 accumulator ( // @[pe.scala 19:29]
    .clock(accumulator_clock),
    .reset(accumulator_reset),
    .io_input_ready(accumulator_io_input_ready),
    .io_input_valid(accumulator_io_input_valid),
    .io_input_bits_x_0(accumulator_io_input_bits_x_0),
    .io_input_bits_last(accumulator_io_input_bits_last),
    .io_output_valid(accumulator_io_output_valid),
    .io_output_bits_x_0(accumulator_io_output_bits_x_0),
    .io_output_bits_last(accumulator_io_output_bits_last)
  );
  Arbiter1ton multiplyOutMux ( // @[pe.scala 20:32]
    .io_input_ready(multiplyOutMux_io_input_ready),
    .io_input_valid(multiplyOutMux_io_input_valid),
    .io_input_bits_x_0(multiplyOutMux_io_input_bits_x_0),
    .io_input_bits_last(multiplyOutMux_io_input_bits_last),
    .io_sel(multiplyOutMux_io_sel),
    .io_output_0_ready(multiplyOutMux_io_output_0_ready),
    .io_output_0_valid(multiplyOutMux_io_output_0_valid),
    .io_output_0_bits_x_0(multiplyOutMux_io_output_0_bits_x_0),
    .io_output_0_bits_last(multiplyOutMux_io_output_0_bits_last),
    .io_output_1_valid(multiplyOutMux_io_output_1_valid),
    .io_output_1_bits_x_0(multiplyOutMux_io_output_1_bits_x_0),
    .io_output_1_bits_last(multiplyOutMux_io_output_1_bits_last)
  );
  Arbiternto1 sumOutMux ( // @[pe.scala 21:27]
    .io_input_0_ready(sumOutMux_io_input_0_ready),
    .io_input_0_valid(sumOutMux_io_input_0_valid),
    .io_input_0_bits_x_0(sumOutMux_io_input_0_bits_x_0),
    .io_input_0_bits_last(sumOutMux_io_input_0_bits_last),
    .io_input_1_valid(sumOutMux_io_input_1_valid),
    .io_input_1_bits_x_0(sumOutMux_io_input_1_bits_x_0),
    .io_input_1_bits_last(sumOutMux_io_input_1_bits_last),
    .io_sel(sumOutMux_io_sel),
    .io_output_ready(sumOutMux_io_output_ready),
    .io_output_valid(sumOutMux_io_output_valid),
    .io_output_bits_x_0(sumOutMux_io_output_bits_x_0),
    .io_output_bits_last(sumOutMux_io_output_bits_last)
  );
  Hsknto1_1 actWeiInHsk ( // @[pecross.scala 14:29]
    .io_input_0_ready(actWeiInHsk_io_input_0_ready),
    .io_input_0_valid(actWeiInHsk_io_input_0_valid),
    .io_input_0_bits_x_0(actWeiInHsk_io_input_0_bits_x_0),
    .io_input_0_bits_last(actWeiInHsk_io_input_0_bits_last),
    .io_input_1_ready(actWeiInHsk_io_input_1_ready),
    .io_input_1_valid(actWeiInHsk_io_input_1_valid),
    .io_input_1_bits_x_0(actWeiInHsk_io_input_1_bits_x_0),
    .io_input_1_bits_last(actWeiInHsk_io_input_1_bits_last),
    .io_output_ready(actWeiInHsk_io_output_ready),
    .io_output_valid(actWeiInHsk_io_output_valid),
    .io_output_bits_0_x_0(actWeiInHsk_io_output_bits_0_x_0),
    .io_output_bits_0_last(actWeiInHsk_io_output_bits_0_last),
    .io_output_bits_1_x_0(actWeiInHsk_io_output_bits_1_x_0),
    .io_output_bits_1_last(actWeiInHsk_io_output_bits_1_last)
  );
  Hsk1ton multiplyInHsk ( // @[pecross.scala 15:31]
    .io_input_ready(multiplyInHsk_io_input_ready),
    .io_input_valid(multiplyInHsk_io_input_valid),
    .io_input_bits_0_x_0(multiplyInHsk_io_input_bits_0_x_0),
    .io_input_bits_0_x_1(multiplyInHsk_io_input_bits_0_x_1),
    .io_input_bits_0_last(multiplyInHsk_io_input_bits_0_last),
    .io_input_bits_1_x_0(multiplyInHsk_io_input_bits_1_x_0),
    .io_input_bits_1_x_1(multiplyInHsk_io_input_bits_1_x_1),
    .io_input_bits_1_last(multiplyInHsk_io_input_bits_1_last),
    .io_input_bits_2_x_0(multiplyInHsk_io_input_bits_2_x_0),
    .io_input_bits_2_x_1(multiplyInHsk_io_input_bits_2_x_1),
    .io_input_bits_2_last(multiplyInHsk_io_input_bits_2_last),
    .io_output_0_ready(multiplyInHsk_io_output_0_ready),
    .io_output_0_valid(multiplyInHsk_io_output_0_valid),
    .io_output_0_bits_x_0(multiplyInHsk_io_output_0_bits_x_0),
    .io_output_0_bits_x_1(multiplyInHsk_io_output_0_bits_x_1),
    .io_output_0_bits_last(multiplyInHsk_io_output_0_bits_last),
    .io_output_1_ready(multiplyInHsk_io_output_1_ready),
    .io_output_1_valid(multiplyInHsk_io_output_1_valid),
    .io_output_1_bits_x_0(multiplyInHsk_io_output_1_bits_x_0),
    .io_output_1_bits_x_1(multiplyInHsk_io_output_1_bits_x_1),
    .io_output_1_bits_last(multiplyInHsk_io_output_1_bits_last),
    .io_output_2_ready(multiplyInHsk_io_output_2_ready),
    .io_output_2_valid(multiplyInHsk_io_output_2_valid),
    .io_output_2_bits_x_0(multiplyInHsk_io_output_2_bits_x_0),
    .io_output_2_bits_x_1(multiplyInHsk_io_output_2_bits_x_1),
    .io_output_2_bits_last(multiplyInHsk_io_output_2_bits_last)
  );
  Arbiternto1_1 weiInMux ( // @[pecross.scala 16:26]
    .io_input_0_ready(weiInMux_io_input_0_ready),
    .io_input_0_valid(weiInMux_io_input_0_valid),
    .io_input_0_bits_x_0(weiInMux_io_input_0_bits_x_0),
    .io_input_0_bits_last(weiInMux_io_input_0_bits_last),
    .io_sel(weiInMux_io_sel),
    .io_output_ready(weiInMux_io_output_ready),
    .io_output_valid(weiInMux_io_output_valid),
    .io_output_bits_x_0(weiInMux_io_output_bits_x_0),
    .io_output_bits_last(weiInMux_io_output_bits_last)
  );
  Arbiternto1_1 actInMux ( // @[pecross.scala 17:26]
    .io_input_0_ready(actInMux_io_input_0_ready),
    .io_input_0_valid(actInMux_io_input_0_valid),
    .io_input_0_bits_x_0(actInMux_io_input_0_bits_x_0),
    .io_input_0_bits_last(actInMux_io_input_0_bits_last),
    .io_sel(actInMux_io_sel),
    .io_output_ready(actInMux_io_output_ready),
    .io_output_valid(actInMux_io_output_valid),
    .io_output_bits_x_0(actInMux_io_output_bits_x_0),
    .io_output_bits_last(actInMux_io_output_bits_last)
  );
  Arbiter1ton_1 multiplyInMux ( // @[pecross.scala 18:31]
    .io_input_ready(multiplyInMux_io_input_ready),
    .io_input_valid(multiplyInMux_io_input_valid),
    .io_input_bits_x_0(multiplyInMux_io_input_bits_x_0),
    .io_input_bits_x_1(multiplyInMux_io_input_bits_x_1),
    .io_input_bits_last(multiplyInMux_io_input_bits_last),
    .io_sel(multiplyInMux_io_sel),
    .io_output_0_ready(multiplyInMux_io_output_0_ready),
    .io_output_0_valid(multiplyInMux_io_output_0_valid),
    .io_output_0_bits_x_0(multiplyInMux_io_output_0_bits_x_0),
    .io_output_0_bits_x_1(multiplyInMux_io_output_0_bits_x_1),
    .io_output_0_bits_last(multiplyInMux_io_output_0_bits_last)
  );
  Arbiter1ton_1 actOutMux ( // @[pecross.scala 19:27]
    .io_input_ready(actOutMux_io_input_ready),
    .io_input_valid(actOutMux_io_input_valid),
    .io_input_bits_x_0(actOutMux_io_input_bits_x_0),
    .io_input_bits_x_1(actOutMux_io_input_bits_x_1),
    .io_input_bits_last(actOutMux_io_input_bits_last),
    .io_sel(actOutMux_io_sel),
    .io_output_0_ready(actOutMux_io_output_0_ready),
    .io_output_0_valid(actOutMux_io_output_0_valid),
    .io_output_0_bits_x_0(actOutMux_io_output_0_bits_x_0),
    .io_output_0_bits_x_1(actOutMux_io_output_0_bits_x_1),
    .io_output_0_bits_last(actOutMux_io_output_0_bits_last)
  );
  Arbiter1ton_1 weiOutMux ( // @[pecross.scala 20:27]
    .io_input_ready(weiOutMux_io_input_ready),
    .io_input_valid(weiOutMux_io_input_valid),
    .io_input_bits_x_0(weiOutMux_io_input_bits_x_0),
    .io_input_bits_x_1(weiOutMux_io_input_bits_x_1),
    .io_input_bits_last(weiOutMux_io_input_bits_last),
    .io_sel(weiOutMux_io_sel),
    .io_output_0_ready(weiOutMux_io_output_0_ready),
    .io_output_0_valid(weiOutMux_io_output_0_valid),
    .io_output_0_bits_x_0(weiOutMux_io_output_0_bits_x_0),
    .io_output_0_bits_x_1(weiOutMux_io_output_0_bits_x_1),
    .io_output_0_bits_last(weiOutMux_io_output_0_bits_last)
  );
  Arbiternto1 adderInMux ( // @[pecross.scala 21:28]
    .io_input_0_ready(adderInMux_io_input_0_ready),
    .io_input_0_valid(adderInMux_io_input_0_valid),
    .io_input_0_bits_x_0(adderInMux_io_input_0_bits_x_0),
    .io_input_0_bits_last(adderInMux_io_input_0_bits_last),
    .io_input_1_valid(adderInMux_io_input_1_valid),
    .io_input_1_bits_x_0(adderInMux_io_input_1_bits_x_0),
    .io_input_1_bits_last(adderInMux_io_input_1_bits_last),
    .io_sel(adderInMux_io_sel),
    .io_output_ready(adderInMux_io_output_ready),
    .io_output_valid(adderInMux_io_output_valid),
    .io_output_bits_x_0(adderInMux_io_output_bits_x_0),
    .io_output_bits_last(adderInMux_io_output_bits_last)
  );
  PipelineHsk actOutHsk ( // @[pecross.scala 47:27]
    .clock(actOutHsk_clock),
    .reset(actOutHsk_reset),
    .io_validPre(actOutHsk_io_validPre),
    .io_readyPre(actOutHsk_io_readyPre),
    .io_lastPre(actOutHsk_io_lastPre),
    .io_validNxt(actOutHsk_io_validNxt),
    .io_readyNxt(actOutHsk_io_readyNxt),
    .io_regen_0(actOutHsk_io_regen_0),
    .io_lastNxt(actOutHsk_io_lastNxt)
  );
  PipelineHsk weiOutHsk ( // @[pecross.scala 58:27]
    .clock(weiOutHsk_clock),
    .reset(weiOutHsk_reset),
    .io_validPre(weiOutHsk_io_validPre),
    .io_readyPre(weiOutHsk_io_readyPre),
    .io_lastPre(weiOutHsk_io_lastPre),
    .io_validNxt(weiOutHsk_io_validNxt),
    .io_readyNxt(weiOutHsk_io_readyNxt),
    .io_regen_0(weiOutHsk_io_regen_0),
    .io_lastNxt(weiOutHsk_io_lastNxt)
  );
  assign multiply_io_input_io_sumIn_ready = adderInHsk_io_input_1_ready; // @[penlr.scala 20:28]
  assign multiply_io_input_io_sumOut_valid = sumOutMux_io_output_valid; // @[pe.scala 29:25]
  assign multiply_io_input_io_sumOut_bits_x_0 = sumOutMux_io_output_bits_x_0; // @[pe.scala 29:25]
  assign multiply_io_input_io_sumOut_bits_last = sumOutMux_io_output_bits_last; // @[pe.scala 29:25]
  assign multiply_io_input_io_actIn_ready = actInMux_io_input_0_ready; // @[pecross.scala 23:14]
  assign multiply_io_input_io_weiIn_ready = weiInMux_io_input_0_ready; // @[pecross.scala 28:14]
  assign multiply_io_input_io_actOut_valid = actOutHsk_io_validNxt; // @[pecross.scala 50:21]
  assign multiply_io_input_io_actOut_bits_x_0 = io_actOut_bits_x_0_r; // @[pecross.scala 54:25]
  assign multiply_io_input_io_actOut_bits_last = actOutHsk_io_lastNxt; // @[pecross.scala 53:25]
  assign multiply_io_input_io_weiOut_valid = weiOutHsk_io_validNxt; // @[pecross.scala 61:21]
  assign multiply_io_input_io_weiOut_bits_x_0 = io_weiOut_bits_x_0_r; // @[pecross.scala 65:25]
  assign multiply_io_input_io_weiOut_bits_last = weiOutHsk_io_lastNxt; // @[pecross.scala 64:25]
  assign multiply_clock = clock;
  assign multiply_reset = reset;
  assign multiply_io_input_valid = multiplyInMux_io_output_0_valid; // @[pecross.scala 42:32]
  assign multiply_io_input_bits_x_0 = multiplyInMux_io_output_0_bits_x_0; // @[pecross.scala 42:32]
  assign multiply_io_input_bits_x_1 = _weiOut_T_1 ? $signed(multiply_io_input_io_weiOut_bits_x_0) : $signed(
    multiplyInMux_io_output_0_bits_x_1); // @[pecross.scala 73:39]
  assign multiply_io_input_bits_last = multiplyInMux_io_output_0_bits_last; // @[pecross.scala 42:32]
  assign multiply_io_output_ready = multiplyOutMux_io_input_ready; // @[pe.scala 24:29]
  assign adder_clock = clock;
  assign adder_reset = reset;
  assign adder_io_input_valid = adderInHsk_io_output_valid; // @[port.scala 24:19]
  assign adder_io_input_bits_x_0 = adderInHsk_io_output_bits_0_x_0; // @[port.scala 20:37]
  assign adder_io_input_bits_x_1 = adderInHsk_io_output_bits_1_x_0; // @[port.scala 20:37]
  assign adder_io_input_bits_last = adderInHsk_io_output_bits_1_last; // @[port.scala 23:23]
  assign adder_io_output_ready = sumOutMux_io_input_0_ready; // @[pe.scala 27:27]
  assign adderInHsk_io_input_0_valid = adderInMux_io_output_valid; // @[pecross.scala 80:26]
  assign adderInHsk_io_input_0_bits_x_0 = adderInMux_io_output_bits_x_0; // @[pecross.scala 80:26]
  assign adderInHsk_io_input_1_valid = multiply_io_input_io_sumIn_valid; // @[penlr.scala 20:28]
  assign adderInHsk_io_input_1_bits_x_0 = multiply_io_input_io_sumIn_bits_x_0; // @[penlr.scala 20:28]
  assign adderInHsk_io_input_1_bits_last = multiply_io_input_io_sumIn_bits_last; // @[penlr.scala 20:28]
  assign adderInHsk_io_output_ready = adder_io_input_ready; // @[port.scala 25:19]
  assign accumulator_clock = clock;
  assign accumulator_reset = reset;
  assign accumulator_io_input_valid = multiplyOutMux_io_output_1_valid; // @[pe.scala 26:33]
  assign accumulator_io_input_bits_x_0 = multiplyOutMux_io_output_1_bits_x_0; // @[pe.scala 26:33]
  assign accumulator_io_input_bits_last = multiplyOutMux_io_output_1_bits_last; // @[pe.scala 26:33]
  assign multiplyOutMux_io_input_valid = multiply_io_output_valid; // @[pe.scala 24:29]
  assign multiplyOutMux_io_input_bits_x_0 = multiply_io_output_bits_x_0; // @[pe.scala 24:29]
  assign multiplyOutMux_io_input_bits_last = multiply_io_output_bits_last; // @[pe.scala 24:29]
  assign multiplyOutMux_io_sel = multiply_io_input_io_statSel == 2'h2 & multiply_io_input_io_actEn; // @[pe.scala 22:53]
  assign multiplyOutMux_io_output_0_ready = adderInMux_io_input_0_ready; // @[pecross.scala 76:33]
  assign sumOutMux_io_input_0_valid = adder_io_output_valid; // @[pe.scala 27:27]
  assign sumOutMux_io_input_0_bits_x_0 = adder_io_output_bits_x_0; // @[pe.scala 27:27]
  assign sumOutMux_io_input_0_bits_last = adder_io_output_bits_last; // @[pe.scala 27:27]
  assign sumOutMux_io_input_1_valid = accumulator_io_output_valid; // @[pe.scala 28:27]
  assign sumOutMux_io_input_1_bits_x_0 = accumulator_io_output_bits_x_0; // @[pe.scala 28:27]
  assign sumOutMux_io_input_1_bits_last = accumulator_io_output_bits_last; // @[pe.scala 28:27]
  assign sumOutMux_io_sel = _multiplyOutMux_io_sel_T & multiply_io_input_io_actEn; // @[pe.scala 23:48]
  assign sumOutMux_io_output_ready = multiply_io_input_io_sumOut_ready; // @[pe.scala 29:25]
  assign actWeiInHsk_io_input_0_valid = actInMux_io_output_valid; // @[pecross.scala 33:24]
  assign actWeiInHsk_io_input_0_bits_x_0 = actInMux_io_output_bits_x_0; // @[pecross.scala 33:24]
  assign actWeiInHsk_io_input_0_bits_last = actInMux_io_output_bits_last; // @[pecross.scala 33:24]
  assign actWeiInHsk_io_input_1_valid = weiInMux_io_output_valid; // @[pecross.scala 34:24]
  assign actWeiInHsk_io_input_1_bits_x_0 = weiInMux_io_output_bits_x_0; // @[pecross.scala 34:24]
  assign actWeiInHsk_io_input_1_bits_last = weiInMux_io_output_bits_last; // @[pecross.scala 34:24]
  assign actWeiInHsk_io_output_ready = multiplyInHsk_io_input_ready; // @[pecross.scala 36:33]
  assign multiplyInHsk_io_input_valid = actWeiInHsk_io_output_valid; // @[pecross.scala 35:34]
  assign multiplyInHsk_io_input_bits_0_x_0 = actWeiInHsk_io_output_bits_0_x_0; // @[port.scala 32:32]
  assign multiplyInHsk_io_input_bits_0_x_1 = actWeiInHsk_io_output_bits_1_x_0; // @[port.scala 32:32]
  assign multiplyInHsk_io_input_bits_0_last = actWeiInHsk_io_output_bits_0_last; // @[port.scala 35:18]
  assign multiplyInHsk_io_input_bits_1_x_0 = actWeiInHsk_io_output_bits_0_x_0; // @[port.scala 32:32]
  assign multiplyInHsk_io_input_bits_1_x_1 = actWeiInHsk_io_output_bits_1_x_0; // @[port.scala 32:32]
  assign multiplyInHsk_io_input_bits_1_last = actWeiInHsk_io_output_bits_0_last; // @[port.scala 35:18]
  assign multiplyInHsk_io_input_bits_2_x_0 = actWeiInHsk_io_output_bits_0_x_0; // @[port.scala 32:32]
  assign multiplyInHsk_io_input_bits_2_x_1 = actWeiInHsk_io_output_bits_1_x_0; // @[port.scala 32:32]
  assign multiplyInHsk_io_input_bits_2_last = actWeiInHsk_io_output_bits_1_last; // @[port.scala 35:18]
  assign multiplyInHsk_io_output_0_ready = multiplyInMux_io_input_ready; // @[pecross.scala 41:28]
  assign multiplyInHsk_io_output_1_ready = actOutMux_io_input_ready; // @[pecross.scala 45:24]
  assign multiplyInHsk_io_output_2_ready = weiOutMux_io_input_ready; // @[pecross.scala 56:24]
  assign weiInMux_io_input_0_valid = multiply_io_input_io_weiIn_valid; // @[pecross.scala 28:14]
  assign weiInMux_io_input_0_bits_x_0 = multiply_io_input_io_weiIn_bits_x_0; // @[pecross.scala 28:14]
  assign weiInMux_io_input_0_bits_last = multiply_io_input_io_weiIn_bits_last; // @[pecross.scala 28:14]
  assign weiInMux_io_sel = _weiOut_T & multiply_io_input_io_weiEn; // @[pecross.scala 69:47]
  assign weiInMux_io_output_ready = actWeiInHsk_io_input_1_ready; // @[pecross.scala 34:24]
  assign actInMux_io_input_0_valid = multiply_io_input_io_actIn_valid; // @[pecross.scala 23:14]
  assign actInMux_io_input_0_bits_x_0 = multiply_io_input_io_actIn_bits_x_0; // @[pecross.scala 23:14]
  assign actInMux_io_input_0_bits_last = multiply_io_input_io_actIn_bits_last; // @[pecross.scala 23:14]
  assign actInMux_io_sel = _weiOut_T & ~multiply_io_input_io_weiEn; // @[pecross.scala 68:47]
  assign actInMux_io_output_ready = actWeiInHsk_io_input_0_ready; // @[pecross.scala 33:24]
  assign multiplyInMux_io_input_valid = multiplyInHsk_io_output_0_valid; // @[pecross.scala 41:28]
  assign multiplyInMux_io_input_bits_x_0 = multiplyInHsk_io_output_0_bits_x_0; // @[pecross.scala 41:28]
  assign multiplyInMux_io_input_bits_x_1 = multiplyInHsk_io_output_0_bits_x_1; // @[pecross.scala 41:28]
  assign multiplyInMux_io_input_bits_last = multiplyInHsk_io_output_0_bits_last; // @[pecross.scala 41:28]
  assign multiplyInMux_io_sel = _weiOut_T & _actInMux_io_sel_T_1; // @[pecross.scala 70:52]
  assign multiplyInMux_io_output_0_ready = multiply_io_input_ready; // @[pecross.scala 42:32]
  assign actOutMux_io_input_valid = multiplyInHsk_io_output_1_valid; // @[pecross.scala 45:24]
  assign actOutMux_io_input_bits_x_0 = multiplyInHsk_io_output_1_bits_x_0; // @[pecross.scala 45:24]
  assign actOutMux_io_input_bits_x_1 = multiplyInHsk_io_output_1_bits_x_1; // @[pecross.scala 45:24]
  assign actOutMux_io_input_bits_last = multiplyInHsk_io_output_1_bits_last; // @[pecross.scala 45:24]
  assign actOutMux_io_sel = _weiOut_T & _actInMux_io_sel_T_1; // @[pecross.scala 71:48]
  assign actOutMux_io_output_0_ready = actOutHsk_io_readyPre; // @[pecross.scala 49:34]
  assign weiOutMux_io_input_valid = multiplyInHsk_io_output_2_valid; // @[pecross.scala 56:24]
  assign weiOutMux_io_input_bits_x_0 = multiplyInHsk_io_output_2_bits_x_0; // @[pecross.scala 56:24]
  assign weiOutMux_io_input_bits_x_1 = multiplyInHsk_io_output_2_bits_x_1; // @[pecross.scala 56:24]
  assign weiOutMux_io_input_bits_last = multiplyInHsk_io_output_2_bits_last; // @[pecross.scala 56:24]
  assign weiOutMux_io_sel = _weiOut_T & multiply_io_input_io_weiEn; // @[pecross.scala 72:48]
  assign weiOutMux_io_output_0_ready = weiOutHsk_io_readyPre; // @[pecross.scala 60:34]
  assign adderInMux_io_input_0_valid = multiplyOutMux_io_output_0_valid; // @[pecross.scala 76:33]
  assign adderInMux_io_input_0_bits_x_0 = multiplyOutMux_io_output_0_bits_x_0; // @[pecross.scala 76:33]
  assign adderInMux_io_input_0_bits_last = multiplyOutMux_io_output_0_bits_last; // @[pecross.scala 76:33]
  assign adderInMux_io_input_1_valid = 1'h1; // @[pecross.scala 77:34]
  assign adderInMux_io_input_1_bits_x_0 = 20'sh0; // @[pecross.scala 78:38]
  assign adderInMux_io_input_1_bits_last = 1'h0; // @[pecross.scala 79:38]
  assign adderInMux_io_sel = _multiplyOutMux_io_sel_T & ~multiply_io_input_io_actEn; // @[pecross.scala 81:49]
  assign adderInMux_io_output_ready = adderInHsk_io_input_0_ready; // @[pecross.scala 80:26]
  assign actOutHsk_clock = clock;
  assign actOutHsk_reset = reset;
  assign actOutHsk_io_validPre = actOutMux_io_output_0_valid; // @[pecross.scala 48:27]
  assign actOutHsk_io_lastPre = actOutMux_io_output_0_bits_last; // @[pecross.scala 52:26]
  assign actOutHsk_io_readyNxt = multiply_io_input_io_actOut_ready; // @[pecross.scala 51:27]
  assign weiOutHsk_clock = clock;
  assign weiOutHsk_reset = reset;
  assign weiOutHsk_io_validPre = weiOutMux_io_output_0_valid; // @[pecross.scala 59:27]
  assign weiOutHsk_io_lastPre = weiOutMux_io_output_0_bits_last; // @[pecross.scala 63:26]
  assign weiOutHsk_io_readyNxt = multiply_io_input_io_weiOut_ready; // @[pecross.scala 62:27]
  always @(posedge clock) begin
    if (actOutHsk_io_regen_0) begin // @[Reg.scala 17:18]
      io_actOut_bits_x_0_r <= actOutMux_io_output_0_bits_x_0; // @[Reg.scala 17:22]
    end
    if (weiOutHsk_io_regen_0) begin // @[Reg.scala 17:18]
      io_weiOut_bits_x_0_r <= weiOutMux_io_output_0_bits_x_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_actOut_bits_x_0_r = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  io_weiOut_bits_x_0_r = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAC(
  input         clock,
  input         reset,
  output        io_actIn_0_ready,
  input         io_actIn_0_valid,
  input  [7:0]  io_actIn_0_bits_x_0,
  input         io_actIn_0_bits_last,
  output        io_actIn_1_ready,
  input         io_actIn_1_valid,
  input  [7:0]  io_actIn_1_bits_x_0,
  input         io_actIn_1_bits_last,
  output        io_actIn_2_ready,
  input         io_actIn_2_valid,
  input  [7:0]  io_actIn_2_bits_x_0,
  input         io_actIn_2_bits_last,
  output        io_actIn_3_ready,
  input         io_actIn_3_valid,
  input  [7:0]  io_actIn_3_bits_x_0,
  input         io_actIn_3_bits_last,
  output        io_actIn_4_ready,
  input         io_actIn_4_valid,
  input  [7:0]  io_actIn_4_bits_x_0,
  input         io_actIn_4_bits_last,
  output        io_actIn_5_ready,
  input         io_actIn_5_valid,
  input  [7:0]  io_actIn_5_bits_x_0,
  input         io_actIn_5_bits_last,
  output        io_actIn_6_ready,
  input         io_actIn_6_valid,
  input  [7:0]  io_actIn_6_bits_x_0,
  input         io_actIn_6_bits_last,
  output        io_actIn_7_ready,
  input         io_actIn_7_valid,
  input  [7:0]  io_actIn_7_bits_x_0,
  input         io_actIn_7_bits_last,
  output        io_actIn_8_ready,
  input         io_actIn_8_valid,
  input  [7:0]  io_actIn_8_bits_x_0,
  input         io_actIn_8_bits_last,
  output        io_actIn_9_ready,
  input         io_actIn_9_valid,
  input  [7:0]  io_actIn_9_bits_x_0,
  input         io_actIn_9_bits_last,
  output        io_actIn_10_ready,
  input         io_actIn_10_valid,
  input  [7:0]  io_actIn_10_bits_x_0,
  input         io_actIn_10_bits_last,
  output        io_actIn_11_ready,
  input         io_actIn_11_valid,
  input  [7:0]  io_actIn_11_bits_x_0,
  input         io_actIn_11_bits_last,
  output        io_actIn_12_ready,
  input         io_actIn_12_valid,
  input  [7:0]  io_actIn_12_bits_x_0,
  input         io_actIn_12_bits_last,
  output        io_actIn_13_ready,
  input         io_actIn_13_valid,
  input  [7:0]  io_actIn_13_bits_x_0,
  input         io_actIn_13_bits_last,
  output        io_actIn_14_ready,
  input         io_actIn_14_valid,
  input  [7:0]  io_actIn_14_bits_x_0,
  input         io_actIn_14_bits_last,
  output        io_actIn_15_ready,
  input         io_actIn_15_valid,
  input  [7:0]  io_actIn_15_bits_x_0,
  input         io_actIn_15_bits_last,
  output        io_weiIn_0_ready,
  input         io_weiIn_0_valid,
  input  [7:0]  io_weiIn_0_bits_x_0,
  input         io_weiIn_0_bits_last,
  output        io_weiIn_1_ready,
  input         io_weiIn_1_valid,
  input  [7:0]  io_weiIn_1_bits_x_0,
  input         io_weiIn_1_bits_last,
  output        io_weiIn_2_ready,
  input         io_weiIn_2_valid,
  input  [7:0]  io_weiIn_2_bits_x_0,
  input         io_weiIn_2_bits_last,
  output        io_weiIn_3_ready,
  input         io_weiIn_3_valid,
  input  [7:0]  io_weiIn_3_bits_x_0,
  input         io_weiIn_3_bits_last,
  output        io_weiIn_4_ready,
  input         io_weiIn_4_valid,
  input  [7:0]  io_weiIn_4_bits_x_0,
  input         io_weiIn_4_bits_last,
  output        io_weiIn_5_ready,
  input         io_weiIn_5_valid,
  input  [7:0]  io_weiIn_5_bits_x_0,
  input         io_weiIn_5_bits_last,
  output        io_weiIn_6_ready,
  input         io_weiIn_6_valid,
  input  [7:0]  io_weiIn_6_bits_x_0,
  input         io_weiIn_6_bits_last,
  output        io_weiIn_7_ready,
  input         io_weiIn_7_valid,
  input  [7:0]  io_weiIn_7_bits_x_0,
  input         io_weiIn_7_bits_last,
  output        io_weiIn_8_ready,
  input         io_weiIn_8_valid,
  input  [7:0]  io_weiIn_8_bits_x_0,
  input         io_weiIn_8_bits_last,
  output        io_weiIn_9_ready,
  input         io_weiIn_9_valid,
  input  [7:0]  io_weiIn_9_bits_x_0,
  input         io_weiIn_9_bits_last,
  output        io_weiIn_10_ready,
  input         io_weiIn_10_valid,
  input  [7:0]  io_weiIn_10_bits_x_0,
  input         io_weiIn_10_bits_last,
  output        io_weiIn_11_ready,
  input         io_weiIn_11_valid,
  input  [7:0]  io_weiIn_11_bits_x_0,
  input         io_weiIn_11_bits_last,
  output        io_weiIn_12_ready,
  input         io_weiIn_12_valid,
  input  [7:0]  io_weiIn_12_bits_x_0,
  input         io_weiIn_12_bits_last,
  output        io_weiIn_13_ready,
  input         io_weiIn_13_valid,
  input  [7:0]  io_weiIn_13_bits_x_0,
  input         io_weiIn_13_bits_last,
  output        io_weiIn_14_ready,
  input         io_weiIn_14_valid,
  input  [7:0]  io_weiIn_14_bits_x_0,
  input         io_weiIn_14_bits_last,
  output        io_weiIn_15_ready,
  input         io_weiIn_15_valid,
  input  [7:0]  io_weiIn_15_bits_x_0,
  input         io_weiIn_15_bits_last,
  output        io_sumIn_0_ready,
  input         io_sumIn_0_valid,
  input  [19:0] io_sumIn_0_bits_x_0,
  input         io_sumIn_0_bits_last,
  output        io_sumIn_1_ready,
  input         io_sumIn_1_valid,
  input  [19:0] io_sumIn_1_bits_x_0,
  input         io_sumIn_1_bits_last,
  output        io_sumIn_2_ready,
  input         io_sumIn_2_valid,
  input  [19:0] io_sumIn_2_bits_x_0,
  input         io_sumIn_2_bits_last,
  output        io_sumIn_3_ready,
  input         io_sumIn_3_valid,
  input  [19:0] io_sumIn_3_bits_x_0,
  input         io_sumIn_3_bits_last,
  output        io_sumIn_4_ready,
  input         io_sumIn_4_valid,
  input  [19:0] io_sumIn_4_bits_x_0,
  input         io_sumIn_4_bits_last,
  output        io_sumIn_5_ready,
  input         io_sumIn_5_valid,
  input  [19:0] io_sumIn_5_bits_x_0,
  input         io_sumIn_5_bits_last,
  output        io_sumIn_6_ready,
  input         io_sumIn_6_valid,
  input  [19:0] io_sumIn_6_bits_x_0,
  input         io_sumIn_6_bits_last,
  output        io_sumIn_7_ready,
  input         io_sumIn_7_valid,
  input  [19:0] io_sumIn_7_bits_x_0,
  input         io_sumIn_7_bits_last,
  output        io_sumIn_8_ready,
  input         io_sumIn_8_valid,
  input  [19:0] io_sumIn_8_bits_x_0,
  input         io_sumIn_8_bits_last,
  output        io_sumIn_9_ready,
  input         io_sumIn_9_valid,
  input  [19:0] io_sumIn_9_bits_x_0,
  input         io_sumIn_9_bits_last,
  output        io_sumIn_10_ready,
  input         io_sumIn_10_valid,
  input  [19:0] io_sumIn_10_bits_x_0,
  input         io_sumIn_10_bits_last,
  output        io_sumIn_11_ready,
  input         io_sumIn_11_valid,
  input  [19:0] io_sumIn_11_bits_x_0,
  input         io_sumIn_11_bits_last,
  output        io_sumIn_12_ready,
  input         io_sumIn_12_valid,
  input  [19:0] io_sumIn_12_bits_x_0,
  input         io_sumIn_12_bits_last,
  output        io_sumIn_13_ready,
  input         io_sumIn_13_valid,
  input  [19:0] io_sumIn_13_bits_x_0,
  input         io_sumIn_13_bits_last,
  output        io_sumIn_14_ready,
  input         io_sumIn_14_valid,
  input  [19:0] io_sumIn_14_bits_x_0,
  input         io_sumIn_14_bits_last,
  output        io_sumIn_15_ready,
  input         io_sumIn_15_valid,
  input  [19:0] io_sumIn_15_bits_x_0,
  input         io_sumIn_15_bits_last,
  input         io_sumOut_0_ready,
  output        io_sumOut_0_valid,
  output [19:0] io_sumOut_0_bits_x_0,
  output        io_sumOut_0_bits_last,
  input         io_sumOut_1_ready,
  output        io_sumOut_1_valid,
  output [19:0] io_sumOut_1_bits_x_0,
  output        io_sumOut_1_bits_last,
  input         io_sumOut_2_ready,
  output        io_sumOut_2_valid,
  output [19:0] io_sumOut_2_bits_x_0,
  output        io_sumOut_2_bits_last,
  input         io_sumOut_3_ready,
  output        io_sumOut_3_valid,
  output [19:0] io_sumOut_3_bits_x_0,
  output        io_sumOut_3_bits_last,
  input         io_sumOut_4_ready,
  output        io_sumOut_4_valid,
  output [19:0] io_sumOut_4_bits_x_0,
  output        io_sumOut_4_bits_last,
  input         io_sumOut_5_ready,
  output        io_sumOut_5_valid,
  output [19:0] io_sumOut_5_bits_x_0,
  output        io_sumOut_5_bits_last,
  input         io_sumOut_6_ready,
  output        io_sumOut_6_valid,
  output [19:0] io_sumOut_6_bits_x_0,
  output        io_sumOut_6_bits_last,
  input         io_sumOut_7_ready,
  output        io_sumOut_7_valid,
  output [19:0] io_sumOut_7_bits_x_0,
  output        io_sumOut_7_bits_last,
  input         io_sumOut_8_ready,
  output        io_sumOut_8_valid,
  output [19:0] io_sumOut_8_bits_x_0,
  output        io_sumOut_8_bits_last,
  input         io_sumOut_9_ready,
  output        io_sumOut_9_valid,
  output [19:0] io_sumOut_9_bits_x_0,
  output        io_sumOut_9_bits_last,
  input         io_sumOut_10_ready,
  output        io_sumOut_10_valid,
  output [19:0] io_sumOut_10_bits_x_0,
  output        io_sumOut_10_bits_last,
  input         io_sumOut_11_ready,
  output        io_sumOut_11_valid,
  output [19:0] io_sumOut_11_bits_x_0,
  output        io_sumOut_11_bits_last,
  input         io_sumOut_12_ready,
  output        io_sumOut_12_valid,
  output [19:0] io_sumOut_12_bits_x_0,
  output        io_sumOut_12_bits_last,
  input         io_sumOut_13_ready,
  output        io_sumOut_13_valid,
  output [19:0] io_sumOut_13_bits_x_0,
  output        io_sumOut_13_bits_last,
  input         io_sumOut_14_ready,
  output        io_sumOut_14_valid,
  output [19:0] io_sumOut_14_bits_x_0,
  output        io_sumOut_14_bits_last,
  input         io_sumOut_15_ready,
  output        io_sumOut_15_valid,
  output [19:0] io_sumOut_15_bits_x_0,
  output        io_sumOut_15_bits_last,
  input  [1:0]  io_statSel,
  input         io_actEn,
  input         io_weiEn,
  input         io_actOutReady,
  input         io_weiOutReady,
  input         rst
);
  wire  PECross_clock; // @[mac.scala 29:63]
  wire  PECross_reset; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_1_clock; // @[mac.scala 29:63]
  wire  PECross_1_reset; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_1_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_1_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_1_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_1_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_1_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_1_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_1_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_1_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_2_clock; // @[mac.scala 29:63]
  wire  PECross_2_reset; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_2_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_2_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_2_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_2_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_2_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_2_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_2_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_2_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_3_clock; // @[mac.scala 29:63]
  wire  PECross_3_reset; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_3_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_3_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_3_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_3_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_3_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_3_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_3_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_3_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_4_clock; // @[mac.scala 29:63]
  wire  PECross_4_reset; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_4_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_4_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_4_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_4_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_4_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_4_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_4_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_4_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_5_clock; // @[mac.scala 29:63]
  wire  PECross_5_reset; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_5_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_5_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_5_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_5_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_5_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_5_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_5_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_5_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_6_clock; // @[mac.scala 29:63]
  wire  PECross_6_reset; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_6_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_6_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_6_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_6_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_6_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_6_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_6_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_6_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_7_clock; // @[mac.scala 29:63]
  wire  PECross_7_reset; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_7_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_7_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_7_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_7_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_7_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_7_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_7_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_7_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_8_clock; // @[mac.scala 29:63]
  wire  PECross_8_reset; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_8_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_8_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_8_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_8_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_8_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_8_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_8_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_8_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_9_clock; // @[mac.scala 29:63]
  wire  PECross_9_reset; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_9_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_9_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_9_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_9_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_9_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_9_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_9_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_9_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_10_clock; // @[mac.scala 29:63]
  wire  PECross_10_reset; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_10_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_10_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_10_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_10_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_10_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_10_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_10_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_10_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_11_clock; // @[mac.scala 29:63]
  wire  PECross_11_reset; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_11_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_11_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_11_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_11_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_11_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_11_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_11_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_11_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_12_clock; // @[mac.scala 29:63]
  wire  PECross_12_reset; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_12_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_12_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_12_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_12_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_12_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_12_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_12_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_12_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_13_clock; // @[mac.scala 29:63]
  wire  PECross_13_reset; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_13_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_13_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_13_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_13_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_13_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_13_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_13_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_13_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_14_clock; // @[mac.scala 29:63]
  wire  PECross_14_reset; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_14_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_14_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_14_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_14_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_14_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_14_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_14_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_14_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_15_clock; // @[mac.scala 29:63]
  wire  PECross_15_reset; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_15_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_15_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_15_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_15_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_15_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_15_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_15_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_15_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_16_clock; // @[mac.scala 29:63]
  wire  PECross_16_reset; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_16_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_16_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_16_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_16_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_16_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_16_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_16_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_16_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_17_clock; // @[mac.scala 29:63]
  wire  PECross_17_reset; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_17_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_17_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_17_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_17_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_17_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_17_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_17_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_17_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_18_clock; // @[mac.scala 29:63]
  wire  PECross_18_reset; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_18_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_18_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_18_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_18_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_18_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_18_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_18_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_18_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_19_clock; // @[mac.scala 29:63]
  wire  PECross_19_reset; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_19_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_19_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_19_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_19_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_19_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_19_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_19_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_19_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_20_clock; // @[mac.scala 29:63]
  wire  PECross_20_reset; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_20_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_20_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_20_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_20_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_20_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_20_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_20_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_20_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_21_clock; // @[mac.scala 29:63]
  wire  PECross_21_reset; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_21_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_21_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_21_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_21_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_21_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_21_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_21_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_21_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_22_clock; // @[mac.scala 29:63]
  wire  PECross_22_reset; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_22_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_22_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_22_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_22_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_22_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_22_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_22_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_22_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_23_clock; // @[mac.scala 29:63]
  wire  PECross_23_reset; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_23_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_23_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_23_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_23_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_23_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_23_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_23_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_23_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_24_clock; // @[mac.scala 29:63]
  wire  PECross_24_reset; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_24_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_24_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_24_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_24_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_24_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_24_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_24_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_24_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_25_clock; // @[mac.scala 29:63]
  wire  PECross_25_reset; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_25_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_25_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_25_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_25_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_25_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_25_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_25_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_25_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_26_clock; // @[mac.scala 29:63]
  wire  PECross_26_reset; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_26_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_26_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_26_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_26_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_26_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_26_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_26_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_26_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_27_clock; // @[mac.scala 29:63]
  wire  PECross_27_reset; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_27_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_27_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_27_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_27_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_27_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_27_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_27_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_27_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_28_clock; // @[mac.scala 29:63]
  wire  PECross_28_reset; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_28_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_28_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_28_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_28_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_28_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_28_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_28_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_28_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_29_clock; // @[mac.scala 29:63]
  wire  PECross_29_reset; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_29_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_29_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_29_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_29_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_29_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_29_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_29_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_29_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_30_clock; // @[mac.scala 29:63]
  wire  PECross_30_reset; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_30_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_30_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_30_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_30_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_30_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_30_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_30_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_30_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_31_clock; // @[mac.scala 29:63]
  wire  PECross_31_reset; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_31_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_31_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_31_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_31_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_31_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_31_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_31_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_31_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_32_clock; // @[mac.scala 29:63]
  wire  PECross_32_reset; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_32_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_32_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_32_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_32_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_32_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_32_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_32_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_32_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_33_clock; // @[mac.scala 29:63]
  wire  PECross_33_reset; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_33_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_33_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_33_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_33_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_33_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_33_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_33_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_33_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_34_clock; // @[mac.scala 29:63]
  wire  PECross_34_reset; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_34_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_34_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_34_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_34_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_34_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_34_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_34_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_34_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_35_clock; // @[mac.scala 29:63]
  wire  PECross_35_reset; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_35_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_35_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_35_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_35_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_35_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_35_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_35_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_35_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_36_clock; // @[mac.scala 29:63]
  wire  PECross_36_reset; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_36_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_36_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_36_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_36_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_36_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_36_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_36_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_36_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_37_clock; // @[mac.scala 29:63]
  wire  PECross_37_reset; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_37_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_37_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_37_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_37_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_37_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_37_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_37_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_37_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_38_clock; // @[mac.scala 29:63]
  wire  PECross_38_reset; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_38_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_38_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_38_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_38_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_38_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_38_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_38_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_38_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_39_clock; // @[mac.scala 29:63]
  wire  PECross_39_reset; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_39_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_39_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_39_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_39_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_39_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_39_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_39_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_39_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_40_clock; // @[mac.scala 29:63]
  wire  PECross_40_reset; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_40_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_40_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_40_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_40_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_40_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_40_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_40_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_40_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_41_clock; // @[mac.scala 29:63]
  wire  PECross_41_reset; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_41_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_41_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_41_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_41_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_41_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_41_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_41_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_41_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_42_clock; // @[mac.scala 29:63]
  wire  PECross_42_reset; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_42_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_42_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_42_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_42_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_42_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_42_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_42_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_42_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_43_clock; // @[mac.scala 29:63]
  wire  PECross_43_reset; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_43_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_43_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_43_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_43_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_43_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_43_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_43_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_43_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_44_clock; // @[mac.scala 29:63]
  wire  PECross_44_reset; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_44_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_44_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_44_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_44_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_44_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_44_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_44_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_44_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_45_clock; // @[mac.scala 29:63]
  wire  PECross_45_reset; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_45_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_45_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_45_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_45_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_45_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_45_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_45_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_45_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_46_clock; // @[mac.scala 29:63]
  wire  PECross_46_reset; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_46_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_46_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_46_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_46_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_46_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_46_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_46_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_46_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_47_clock; // @[mac.scala 29:63]
  wire  PECross_47_reset; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_47_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_47_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_47_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_47_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_47_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_47_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_47_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_47_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_48_clock; // @[mac.scala 29:63]
  wire  PECross_48_reset; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_48_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_48_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_48_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_48_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_48_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_48_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_48_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_48_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_49_clock; // @[mac.scala 29:63]
  wire  PECross_49_reset; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_49_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_49_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_49_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_49_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_49_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_49_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_49_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_49_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_50_clock; // @[mac.scala 29:63]
  wire  PECross_50_reset; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_50_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_50_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_50_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_50_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_50_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_50_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_50_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_50_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_51_clock; // @[mac.scala 29:63]
  wire  PECross_51_reset; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_51_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_51_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_51_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_51_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_51_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_51_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_51_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_51_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_52_clock; // @[mac.scala 29:63]
  wire  PECross_52_reset; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_52_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_52_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_52_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_52_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_52_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_52_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_52_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_52_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_53_clock; // @[mac.scala 29:63]
  wire  PECross_53_reset; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_53_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_53_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_53_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_53_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_53_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_53_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_53_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_53_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_54_clock; // @[mac.scala 29:63]
  wire  PECross_54_reset; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_54_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_54_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_54_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_54_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_54_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_54_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_54_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_54_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_55_clock; // @[mac.scala 29:63]
  wire  PECross_55_reset; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_55_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_55_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_55_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_55_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_55_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_55_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_55_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_55_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_56_clock; // @[mac.scala 29:63]
  wire  PECross_56_reset; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_56_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_56_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_56_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_56_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_56_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_56_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_56_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_56_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_57_clock; // @[mac.scala 29:63]
  wire  PECross_57_reset; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_57_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_57_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_57_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_57_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_57_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_57_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_57_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_57_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_58_clock; // @[mac.scala 29:63]
  wire  PECross_58_reset; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_58_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_58_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_58_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_58_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_58_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_58_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_58_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_58_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_59_clock; // @[mac.scala 29:63]
  wire  PECross_59_reset; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_59_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_59_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_59_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_59_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_59_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_59_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_59_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_59_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_60_clock; // @[mac.scala 29:63]
  wire  PECross_60_reset; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_60_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_60_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_60_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_60_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_60_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_60_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_60_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_60_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_61_clock; // @[mac.scala 29:63]
  wire  PECross_61_reset; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_61_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_61_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_61_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_61_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_61_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_61_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_61_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_61_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_62_clock; // @[mac.scala 29:63]
  wire  PECross_62_reset; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_62_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_62_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_62_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_62_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_62_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_62_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_62_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_62_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_63_clock; // @[mac.scala 29:63]
  wire  PECross_63_reset; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_63_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_63_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_63_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_63_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_63_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_63_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_63_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_63_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_64_clock; // @[mac.scala 29:63]
  wire  PECross_64_reset; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_64_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_64_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_64_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_64_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_64_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_64_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_64_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_64_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_65_clock; // @[mac.scala 29:63]
  wire  PECross_65_reset; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_65_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_65_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_65_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_65_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_65_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_65_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_65_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_65_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_66_clock; // @[mac.scala 29:63]
  wire  PECross_66_reset; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_66_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_66_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_66_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_66_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_66_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_66_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_66_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_66_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_67_clock; // @[mac.scala 29:63]
  wire  PECross_67_reset; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_67_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_67_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_67_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_67_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_67_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_67_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_67_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_67_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_68_clock; // @[mac.scala 29:63]
  wire  PECross_68_reset; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_68_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_68_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_68_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_68_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_68_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_68_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_68_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_68_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_69_clock; // @[mac.scala 29:63]
  wire  PECross_69_reset; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_69_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_69_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_69_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_69_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_69_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_69_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_69_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_69_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_70_clock; // @[mac.scala 29:63]
  wire  PECross_70_reset; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_70_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_70_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_70_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_70_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_70_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_70_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_70_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_70_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_71_clock; // @[mac.scala 29:63]
  wire  PECross_71_reset; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_71_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_71_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_71_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_71_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_71_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_71_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_71_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_71_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_72_clock; // @[mac.scala 29:63]
  wire  PECross_72_reset; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_72_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_72_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_72_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_72_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_72_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_72_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_72_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_72_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_73_clock; // @[mac.scala 29:63]
  wire  PECross_73_reset; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_73_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_73_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_73_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_73_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_73_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_73_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_73_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_73_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_74_clock; // @[mac.scala 29:63]
  wire  PECross_74_reset; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_74_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_74_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_74_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_74_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_74_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_74_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_74_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_74_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_75_clock; // @[mac.scala 29:63]
  wire  PECross_75_reset; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_75_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_75_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_75_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_75_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_75_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_75_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_75_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_75_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_76_clock; // @[mac.scala 29:63]
  wire  PECross_76_reset; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_76_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_76_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_76_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_76_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_76_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_76_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_76_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_76_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_77_clock; // @[mac.scala 29:63]
  wire  PECross_77_reset; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_77_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_77_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_77_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_77_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_77_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_77_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_77_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_77_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_78_clock; // @[mac.scala 29:63]
  wire  PECross_78_reset; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_78_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_78_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_78_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_78_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_78_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_78_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_78_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_78_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_79_clock; // @[mac.scala 29:63]
  wire  PECross_79_reset; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_79_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_79_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_79_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_79_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_79_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_79_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_79_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_79_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_80_clock; // @[mac.scala 29:63]
  wire  PECross_80_reset; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_80_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_80_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_80_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_80_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_80_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_80_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_80_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_80_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_81_clock; // @[mac.scala 29:63]
  wire  PECross_81_reset; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_81_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_81_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_81_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_81_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_81_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_81_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_81_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_81_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_82_clock; // @[mac.scala 29:63]
  wire  PECross_82_reset; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_82_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_82_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_82_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_82_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_82_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_82_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_82_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_82_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_83_clock; // @[mac.scala 29:63]
  wire  PECross_83_reset; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_83_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_83_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_83_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_83_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_83_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_83_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_83_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_83_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_84_clock; // @[mac.scala 29:63]
  wire  PECross_84_reset; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_84_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_84_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_84_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_84_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_84_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_84_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_84_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_84_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_85_clock; // @[mac.scala 29:63]
  wire  PECross_85_reset; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_85_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_85_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_85_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_85_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_85_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_85_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_85_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_85_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_86_clock; // @[mac.scala 29:63]
  wire  PECross_86_reset; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_86_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_86_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_86_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_86_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_86_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_86_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_86_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_86_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_87_clock; // @[mac.scala 29:63]
  wire  PECross_87_reset; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_87_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_87_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_87_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_87_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_87_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_87_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_87_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_87_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_88_clock; // @[mac.scala 29:63]
  wire  PECross_88_reset; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_88_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_88_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_88_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_88_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_88_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_88_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_88_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_88_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_89_clock; // @[mac.scala 29:63]
  wire  PECross_89_reset; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_89_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_89_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_89_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_89_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_89_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_89_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_89_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_89_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_90_clock; // @[mac.scala 29:63]
  wire  PECross_90_reset; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_90_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_90_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_90_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_90_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_90_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_90_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_90_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_90_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_91_clock; // @[mac.scala 29:63]
  wire  PECross_91_reset; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_91_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_91_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_91_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_91_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_91_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_91_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_91_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_91_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_92_clock; // @[mac.scala 29:63]
  wire  PECross_92_reset; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_92_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_92_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_92_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_92_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_92_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_92_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_92_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_92_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_93_clock; // @[mac.scala 29:63]
  wire  PECross_93_reset; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_93_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_93_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_93_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_93_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_93_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_93_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_93_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_93_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_94_clock; // @[mac.scala 29:63]
  wire  PECross_94_reset; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_94_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_94_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_94_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_94_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_94_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_94_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_94_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_94_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_95_clock; // @[mac.scala 29:63]
  wire  PECross_95_reset; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_95_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_95_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_95_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_95_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_95_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_95_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_95_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_95_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_96_clock; // @[mac.scala 29:63]
  wire  PECross_96_reset; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_96_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_96_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_96_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_96_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_96_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_96_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_96_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_96_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_97_clock; // @[mac.scala 29:63]
  wire  PECross_97_reset; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_97_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_97_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_97_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_97_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_97_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_97_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_97_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_97_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_98_clock; // @[mac.scala 29:63]
  wire  PECross_98_reset; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_98_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_98_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_98_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_98_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_98_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_98_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_98_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_98_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_99_clock; // @[mac.scala 29:63]
  wire  PECross_99_reset; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_99_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_99_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_99_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_99_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_99_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_99_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_99_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_99_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_100_clock; // @[mac.scala 29:63]
  wire  PECross_100_reset; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_100_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_100_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_100_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_100_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_100_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_100_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_100_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_100_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_101_clock; // @[mac.scala 29:63]
  wire  PECross_101_reset; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_101_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_101_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_101_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_101_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_101_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_101_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_101_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_101_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_102_clock; // @[mac.scala 29:63]
  wire  PECross_102_reset; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_102_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_102_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_102_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_102_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_102_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_102_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_102_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_102_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_103_clock; // @[mac.scala 29:63]
  wire  PECross_103_reset; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_103_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_103_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_103_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_103_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_103_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_103_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_103_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_103_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_104_clock; // @[mac.scala 29:63]
  wire  PECross_104_reset; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_104_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_104_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_104_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_104_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_104_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_104_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_104_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_104_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_105_clock; // @[mac.scala 29:63]
  wire  PECross_105_reset; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_105_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_105_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_105_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_105_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_105_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_105_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_105_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_105_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_106_clock; // @[mac.scala 29:63]
  wire  PECross_106_reset; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_106_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_106_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_106_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_106_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_106_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_106_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_106_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_106_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_107_clock; // @[mac.scala 29:63]
  wire  PECross_107_reset; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_107_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_107_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_107_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_107_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_107_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_107_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_107_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_107_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_108_clock; // @[mac.scala 29:63]
  wire  PECross_108_reset; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_108_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_108_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_108_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_108_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_108_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_108_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_108_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_108_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_109_clock; // @[mac.scala 29:63]
  wire  PECross_109_reset; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_109_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_109_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_109_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_109_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_109_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_109_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_109_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_109_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_110_clock; // @[mac.scala 29:63]
  wire  PECross_110_reset; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_110_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_110_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_110_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_110_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_110_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_110_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_110_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_110_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_111_clock; // @[mac.scala 29:63]
  wire  PECross_111_reset; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_111_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_111_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_111_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_111_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_111_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_111_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_111_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_111_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_112_clock; // @[mac.scala 29:63]
  wire  PECross_112_reset; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_112_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_112_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_112_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_112_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_112_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_112_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_112_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_112_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_113_clock; // @[mac.scala 29:63]
  wire  PECross_113_reset; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_113_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_113_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_113_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_113_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_113_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_113_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_113_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_113_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_114_clock; // @[mac.scala 29:63]
  wire  PECross_114_reset; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_114_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_114_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_114_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_114_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_114_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_114_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_114_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_114_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_115_clock; // @[mac.scala 29:63]
  wire  PECross_115_reset; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_115_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_115_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_115_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_115_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_115_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_115_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_115_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_115_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_116_clock; // @[mac.scala 29:63]
  wire  PECross_116_reset; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_116_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_116_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_116_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_116_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_116_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_116_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_116_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_116_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_117_clock; // @[mac.scala 29:63]
  wire  PECross_117_reset; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_117_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_117_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_117_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_117_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_117_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_117_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_117_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_117_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_118_clock; // @[mac.scala 29:63]
  wire  PECross_118_reset; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_118_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_118_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_118_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_118_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_118_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_118_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_118_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_118_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_119_clock; // @[mac.scala 29:63]
  wire  PECross_119_reset; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_119_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_119_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_119_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_119_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_119_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_119_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_119_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_119_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_120_clock; // @[mac.scala 29:63]
  wire  PECross_120_reset; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_120_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_120_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_120_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_120_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_120_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_120_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_120_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_120_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_121_clock; // @[mac.scala 29:63]
  wire  PECross_121_reset; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_121_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_121_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_121_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_121_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_121_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_121_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_121_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_121_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_122_clock; // @[mac.scala 29:63]
  wire  PECross_122_reset; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_122_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_122_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_122_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_122_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_122_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_122_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_122_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_122_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_123_clock; // @[mac.scala 29:63]
  wire  PECross_123_reset; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_123_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_123_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_123_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_123_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_123_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_123_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_123_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_123_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_124_clock; // @[mac.scala 29:63]
  wire  PECross_124_reset; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_124_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_124_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_124_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_124_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_124_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_124_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_124_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_124_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_125_clock; // @[mac.scala 29:63]
  wire  PECross_125_reset; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_125_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_125_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_125_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_125_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_125_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_125_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_125_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_125_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_126_clock; // @[mac.scala 29:63]
  wire  PECross_126_reset; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_126_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_126_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_126_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_126_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_126_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_126_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_126_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_126_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_127_clock; // @[mac.scala 29:63]
  wire  PECross_127_reset; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_127_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_127_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_127_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_127_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_127_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_127_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_127_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_127_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_128_clock; // @[mac.scala 29:63]
  wire  PECross_128_reset; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_128_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_128_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_128_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_128_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_128_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_128_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_128_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_128_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_129_clock; // @[mac.scala 29:63]
  wire  PECross_129_reset; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_129_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_129_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_129_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_129_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_129_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_129_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_129_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_129_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_130_clock; // @[mac.scala 29:63]
  wire  PECross_130_reset; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_130_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_130_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_130_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_130_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_130_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_130_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_130_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_130_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_131_clock; // @[mac.scala 29:63]
  wire  PECross_131_reset; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_131_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_131_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_131_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_131_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_131_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_131_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_131_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_131_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_132_clock; // @[mac.scala 29:63]
  wire  PECross_132_reset; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_132_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_132_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_132_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_132_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_132_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_132_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_132_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_132_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_133_clock; // @[mac.scala 29:63]
  wire  PECross_133_reset; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_133_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_133_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_133_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_133_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_133_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_133_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_133_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_133_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_134_clock; // @[mac.scala 29:63]
  wire  PECross_134_reset; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_134_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_134_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_134_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_134_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_134_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_134_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_134_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_134_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_135_clock; // @[mac.scala 29:63]
  wire  PECross_135_reset; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_135_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_135_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_135_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_135_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_135_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_135_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_135_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_135_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_136_clock; // @[mac.scala 29:63]
  wire  PECross_136_reset; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_136_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_136_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_136_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_136_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_136_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_136_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_136_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_136_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_137_clock; // @[mac.scala 29:63]
  wire  PECross_137_reset; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_137_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_137_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_137_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_137_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_137_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_137_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_137_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_137_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_138_clock; // @[mac.scala 29:63]
  wire  PECross_138_reset; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_138_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_138_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_138_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_138_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_138_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_138_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_138_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_138_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_139_clock; // @[mac.scala 29:63]
  wire  PECross_139_reset; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_139_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_139_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_139_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_139_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_139_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_139_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_139_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_139_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_140_clock; // @[mac.scala 29:63]
  wire  PECross_140_reset; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_140_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_140_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_140_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_140_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_140_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_140_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_140_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_140_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_141_clock; // @[mac.scala 29:63]
  wire  PECross_141_reset; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_141_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_141_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_141_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_141_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_141_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_141_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_141_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_141_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_142_clock; // @[mac.scala 29:63]
  wire  PECross_142_reset; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_142_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_142_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_142_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_142_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_142_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_142_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_142_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_142_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_143_clock; // @[mac.scala 29:63]
  wire  PECross_143_reset; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_143_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_143_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_143_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_143_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_143_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_143_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_143_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_143_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_144_clock; // @[mac.scala 29:63]
  wire  PECross_144_reset; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_144_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_144_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_144_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_144_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_144_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_144_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_144_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_144_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_145_clock; // @[mac.scala 29:63]
  wire  PECross_145_reset; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_145_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_145_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_145_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_145_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_145_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_145_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_145_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_145_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_146_clock; // @[mac.scala 29:63]
  wire  PECross_146_reset; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_146_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_146_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_146_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_146_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_146_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_146_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_146_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_146_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_147_clock; // @[mac.scala 29:63]
  wire  PECross_147_reset; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_147_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_147_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_147_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_147_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_147_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_147_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_147_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_147_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_148_clock; // @[mac.scala 29:63]
  wire  PECross_148_reset; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_148_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_148_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_148_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_148_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_148_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_148_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_148_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_148_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_149_clock; // @[mac.scala 29:63]
  wire  PECross_149_reset; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_149_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_149_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_149_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_149_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_149_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_149_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_149_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_149_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_150_clock; // @[mac.scala 29:63]
  wire  PECross_150_reset; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_150_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_150_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_150_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_150_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_150_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_150_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_150_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_150_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_151_clock; // @[mac.scala 29:63]
  wire  PECross_151_reset; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_151_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_151_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_151_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_151_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_151_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_151_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_151_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_151_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_152_clock; // @[mac.scala 29:63]
  wire  PECross_152_reset; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_152_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_152_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_152_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_152_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_152_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_152_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_152_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_152_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_153_clock; // @[mac.scala 29:63]
  wire  PECross_153_reset; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_153_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_153_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_153_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_153_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_153_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_153_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_153_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_153_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_154_clock; // @[mac.scala 29:63]
  wire  PECross_154_reset; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_154_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_154_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_154_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_154_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_154_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_154_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_154_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_154_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_155_clock; // @[mac.scala 29:63]
  wire  PECross_155_reset; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_155_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_155_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_155_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_155_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_155_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_155_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_155_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_155_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_156_clock; // @[mac.scala 29:63]
  wire  PECross_156_reset; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_156_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_156_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_156_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_156_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_156_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_156_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_156_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_156_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_157_clock; // @[mac.scala 29:63]
  wire  PECross_157_reset; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_157_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_157_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_157_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_157_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_157_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_157_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_157_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_157_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_158_clock; // @[mac.scala 29:63]
  wire  PECross_158_reset; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_158_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_158_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_158_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_158_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_158_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_158_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_158_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_158_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_159_clock; // @[mac.scala 29:63]
  wire  PECross_159_reset; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_159_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_159_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_159_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_159_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_159_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_159_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_159_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_159_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_160_clock; // @[mac.scala 29:63]
  wire  PECross_160_reset; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_160_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_160_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_160_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_160_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_160_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_160_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_160_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_160_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_161_clock; // @[mac.scala 29:63]
  wire  PECross_161_reset; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_161_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_161_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_161_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_161_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_161_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_161_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_161_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_161_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_162_clock; // @[mac.scala 29:63]
  wire  PECross_162_reset; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_162_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_162_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_162_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_162_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_162_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_162_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_162_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_162_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_163_clock; // @[mac.scala 29:63]
  wire  PECross_163_reset; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_163_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_163_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_163_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_163_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_163_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_163_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_163_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_163_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_164_clock; // @[mac.scala 29:63]
  wire  PECross_164_reset; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_164_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_164_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_164_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_164_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_164_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_164_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_164_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_164_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_165_clock; // @[mac.scala 29:63]
  wire  PECross_165_reset; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_165_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_165_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_165_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_165_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_165_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_165_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_165_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_165_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_166_clock; // @[mac.scala 29:63]
  wire  PECross_166_reset; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_166_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_166_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_166_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_166_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_166_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_166_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_166_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_166_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_167_clock; // @[mac.scala 29:63]
  wire  PECross_167_reset; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_167_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_167_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_167_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_167_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_167_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_167_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_167_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_167_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_168_clock; // @[mac.scala 29:63]
  wire  PECross_168_reset; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_168_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_168_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_168_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_168_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_168_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_168_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_168_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_168_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_169_clock; // @[mac.scala 29:63]
  wire  PECross_169_reset; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_169_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_169_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_169_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_169_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_169_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_169_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_169_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_169_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_170_clock; // @[mac.scala 29:63]
  wire  PECross_170_reset; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_170_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_170_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_170_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_170_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_170_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_170_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_170_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_170_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_171_clock; // @[mac.scala 29:63]
  wire  PECross_171_reset; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_171_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_171_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_171_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_171_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_171_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_171_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_171_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_171_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_172_clock; // @[mac.scala 29:63]
  wire  PECross_172_reset; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_172_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_172_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_172_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_172_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_172_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_172_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_172_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_172_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_173_clock; // @[mac.scala 29:63]
  wire  PECross_173_reset; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_173_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_173_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_173_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_173_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_173_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_173_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_173_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_173_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_174_clock; // @[mac.scala 29:63]
  wire  PECross_174_reset; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_174_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_174_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_174_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_174_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_174_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_174_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_174_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_174_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_175_clock; // @[mac.scala 29:63]
  wire  PECross_175_reset; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_175_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_175_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_175_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_175_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_175_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_175_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_175_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_175_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_176_clock; // @[mac.scala 29:63]
  wire  PECross_176_reset; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_176_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_176_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_176_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_176_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_176_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_176_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_176_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_176_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_177_clock; // @[mac.scala 29:63]
  wire  PECross_177_reset; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_177_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_177_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_177_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_177_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_177_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_177_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_177_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_177_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_178_clock; // @[mac.scala 29:63]
  wire  PECross_178_reset; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_178_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_178_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_178_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_178_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_178_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_178_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_178_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_178_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_179_clock; // @[mac.scala 29:63]
  wire  PECross_179_reset; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_179_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_179_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_179_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_179_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_179_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_179_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_179_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_179_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_180_clock; // @[mac.scala 29:63]
  wire  PECross_180_reset; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_180_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_180_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_180_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_180_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_180_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_180_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_180_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_180_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_181_clock; // @[mac.scala 29:63]
  wire  PECross_181_reset; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_181_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_181_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_181_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_181_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_181_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_181_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_181_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_181_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_182_clock; // @[mac.scala 29:63]
  wire  PECross_182_reset; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_182_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_182_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_182_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_182_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_182_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_182_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_182_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_182_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_183_clock; // @[mac.scala 29:63]
  wire  PECross_183_reset; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_183_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_183_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_183_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_183_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_183_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_183_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_183_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_183_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_184_clock; // @[mac.scala 29:63]
  wire  PECross_184_reset; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_184_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_184_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_184_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_184_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_184_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_184_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_184_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_184_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_185_clock; // @[mac.scala 29:63]
  wire  PECross_185_reset; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_185_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_185_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_185_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_185_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_185_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_185_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_185_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_185_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_186_clock; // @[mac.scala 29:63]
  wire  PECross_186_reset; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_186_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_186_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_186_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_186_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_186_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_186_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_186_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_186_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_187_clock; // @[mac.scala 29:63]
  wire  PECross_187_reset; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_187_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_187_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_187_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_187_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_187_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_187_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_187_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_187_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_188_clock; // @[mac.scala 29:63]
  wire  PECross_188_reset; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_188_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_188_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_188_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_188_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_188_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_188_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_188_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_188_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_189_clock; // @[mac.scala 29:63]
  wire  PECross_189_reset; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_189_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_189_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_189_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_189_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_189_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_189_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_189_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_189_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_190_clock; // @[mac.scala 29:63]
  wire  PECross_190_reset; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_190_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_190_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_190_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_190_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_190_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_190_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_190_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_190_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_191_clock; // @[mac.scala 29:63]
  wire  PECross_191_reset; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_191_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_191_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_191_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_191_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_191_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_191_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_191_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_191_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_192_clock; // @[mac.scala 29:63]
  wire  PECross_192_reset; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_192_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_192_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_192_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_192_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_192_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_192_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_192_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_192_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_193_clock; // @[mac.scala 29:63]
  wire  PECross_193_reset; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_193_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_193_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_193_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_193_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_193_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_193_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_193_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_193_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_194_clock; // @[mac.scala 29:63]
  wire  PECross_194_reset; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_194_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_194_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_194_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_194_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_194_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_194_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_194_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_194_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_195_clock; // @[mac.scala 29:63]
  wire  PECross_195_reset; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_195_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_195_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_195_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_195_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_195_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_195_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_195_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_195_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_196_clock; // @[mac.scala 29:63]
  wire  PECross_196_reset; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_196_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_196_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_196_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_196_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_196_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_196_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_196_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_196_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_197_clock; // @[mac.scala 29:63]
  wire  PECross_197_reset; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_197_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_197_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_197_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_197_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_197_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_197_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_197_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_197_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_198_clock; // @[mac.scala 29:63]
  wire  PECross_198_reset; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_198_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_198_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_198_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_198_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_198_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_198_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_198_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_198_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_199_clock; // @[mac.scala 29:63]
  wire  PECross_199_reset; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_199_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_199_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_199_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_199_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_199_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_199_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_199_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_199_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_200_clock; // @[mac.scala 29:63]
  wire  PECross_200_reset; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_200_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_200_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_200_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_200_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_200_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_200_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_200_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_200_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_201_clock; // @[mac.scala 29:63]
  wire  PECross_201_reset; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_201_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_201_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_201_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_201_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_201_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_201_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_201_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_201_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_202_clock; // @[mac.scala 29:63]
  wire  PECross_202_reset; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_202_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_202_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_202_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_202_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_202_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_202_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_202_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_202_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_203_clock; // @[mac.scala 29:63]
  wire  PECross_203_reset; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_203_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_203_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_203_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_203_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_203_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_203_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_203_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_203_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_204_clock; // @[mac.scala 29:63]
  wire  PECross_204_reset; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_204_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_204_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_204_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_204_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_204_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_204_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_204_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_204_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_205_clock; // @[mac.scala 29:63]
  wire  PECross_205_reset; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_205_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_205_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_205_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_205_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_205_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_205_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_205_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_205_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_206_clock; // @[mac.scala 29:63]
  wire  PECross_206_reset; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_206_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_206_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_206_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_206_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_206_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_206_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_206_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_206_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_207_clock; // @[mac.scala 29:63]
  wire  PECross_207_reset; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_207_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_207_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_207_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_207_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_207_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_207_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_207_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_207_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_208_clock; // @[mac.scala 29:63]
  wire  PECross_208_reset; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_208_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_208_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_208_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_208_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_208_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_208_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_208_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_208_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_209_clock; // @[mac.scala 29:63]
  wire  PECross_209_reset; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_209_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_209_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_209_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_209_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_209_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_209_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_209_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_209_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_210_clock; // @[mac.scala 29:63]
  wire  PECross_210_reset; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_210_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_210_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_210_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_210_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_210_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_210_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_210_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_210_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_211_clock; // @[mac.scala 29:63]
  wire  PECross_211_reset; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_211_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_211_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_211_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_211_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_211_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_211_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_211_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_211_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_212_clock; // @[mac.scala 29:63]
  wire  PECross_212_reset; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_212_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_212_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_212_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_212_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_212_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_212_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_212_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_212_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_213_clock; // @[mac.scala 29:63]
  wire  PECross_213_reset; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_213_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_213_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_213_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_213_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_213_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_213_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_213_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_213_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_214_clock; // @[mac.scala 29:63]
  wire  PECross_214_reset; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_214_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_214_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_214_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_214_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_214_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_214_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_214_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_214_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_215_clock; // @[mac.scala 29:63]
  wire  PECross_215_reset; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_215_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_215_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_215_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_215_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_215_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_215_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_215_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_215_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_216_clock; // @[mac.scala 29:63]
  wire  PECross_216_reset; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_216_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_216_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_216_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_216_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_216_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_216_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_216_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_216_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_217_clock; // @[mac.scala 29:63]
  wire  PECross_217_reset; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_217_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_217_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_217_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_217_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_217_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_217_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_217_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_217_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_218_clock; // @[mac.scala 29:63]
  wire  PECross_218_reset; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_218_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_218_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_218_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_218_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_218_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_218_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_218_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_218_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_219_clock; // @[mac.scala 29:63]
  wire  PECross_219_reset; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_219_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_219_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_219_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_219_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_219_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_219_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_219_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_219_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_220_clock; // @[mac.scala 29:63]
  wire  PECross_220_reset; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_220_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_220_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_220_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_220_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_220_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_220_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_220_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_220_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_221_clock; // @[mac.scala 29:63]
  wire  PECross_221_reset; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_221_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_221_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_221_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_221_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_221_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_221_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_221_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_221_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_222_clock; // @[mac.scala 29:63]
  wire  PECross_222_reset; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_222_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_222_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_222_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_222_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_222_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_222_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_222_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_222_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_223_clock; // @[mac.scala 29:63]
  wire  PECross_223_reset; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_223_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_223_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_223_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_223_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_223_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_223_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_223_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_223_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_224_clock; // @[mac.scala 29:63]
  wire  PECross_224_reset; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_224_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_224_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_224_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_224_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_224_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_224_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_224_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_224_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_225_clock; // @[mac.scala 29:63]
  wire  PECross_225_reset; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_225_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_225_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_225_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_225_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_225_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_225_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_225_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_225_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_226_clock; // @[mac.scala 29:63]
  wire  PECross_226_reset; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_226_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_226_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_226_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_226_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_226_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_226_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_226_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_226_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_227_clock; // @[mac.scala 29:63]
  wire  PECross_227_reset; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_227_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_227_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_227_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_227_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_227_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_227_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_227_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_227_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_228_clock; // @[mac.scala 29:63]
  wire  PECross_228_reset; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_228_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_228_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_228_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_228_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_228_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_228_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_228_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_228_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_229_clock; // @[mac.scala 29:63]
  wire  PECross_229_reset; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_229_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_229_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_229_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_229_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_229_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_229_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_229_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_229_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_230_clock; // @[mac.scala 29:63]
  wire  PECross_230_reset; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_230_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_230_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_230_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_230_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_230_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_230_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_230_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_230_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_231_clock; // @[mac.scala 29:63]
  wire  PECross_231_reset; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_231_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_231_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_231_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_231_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_231_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_231_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_231_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_231_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_232_clock; // @[mac.scala 29:63]
  wire  PECross_232_reset; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_232_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_232_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_232_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_232_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_232_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_232_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_232_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_232_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_233_clock; // @[mac.scala 29:63]
  wire  PECross_233_reset; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_233_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_233_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_233_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_233_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_233_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_233_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_233_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_233_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_234_clock; // @[mac.scala 29:63]
  wire  PECross_234_reset; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_234_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_234_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_234_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_234_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_234_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_234_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_234_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_234_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_235_clock; // @[mac.scala 29:63]
  wire  PECross_235_reset; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_235_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_235_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_235_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_235_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_235_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_235_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_235_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_235_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_236_clock; // @[mac.scala 29:63]
  wire  PECross_236_reset; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_236_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_236_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_236_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_236_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_236_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_236_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_236_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_236_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_237_clock; // @[mac.scala 29:63]
  wire  PECross_237_reset; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_237_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_237_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_237_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_237_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_237_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_237_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_237_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_237_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_238_clock; // @[mac.scala 29:63]
  wire  PECross_238_reset; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_238_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_238_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_238_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_238_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_238_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_238_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_238_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_238_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_239_clock; // @[mac.scala 29:63]
  wire  PECross_239_reset; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_239_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_239_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_239_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_239_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_239_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_239_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_239_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_239_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_240_clock; // @[mac.scala 29:63]
  wire  PECross_240_reset; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_240_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_240_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_240_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_240_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_240_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_240_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_240_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_240_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_241_clock; // @[mac.scala 29:63]
  wire  PECross_241_reset; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_241_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_241_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_241_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_241_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_241_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_241_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_241_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_241_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_242_clock; // @[mac.scala 29:63]
  wire  PECross_242_reset; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_242_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_242_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_242_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_242_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_242_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_242_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_242_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_242_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_243_clock; // @[mac.scala 29:63]
  wire  PECross_243_reset; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_243_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_243_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_243_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_243_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_243_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_243_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_243_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_243_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_244_clock; // @[mac.scala 29:63]
  wire  PECross_244_reset; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_244_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_244_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_244_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_244_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_244_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_244_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_244_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_244_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_245_clock; // @[mac.scala 29:63]
  wire  PECross_245_reset; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_245_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_245_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_245_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_245_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_245_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_245_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_245_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_245_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_246_clock; // @[mac.scala 29:63]
  wire  PECross_246_reset; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_246_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_246_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_246_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_246_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_246_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_246_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_246_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_246_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_247_clock; // @[mac.scala 29:63]
  wire  PECross_247_reset; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_247_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_247_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_247_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_247_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_247_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_247_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_247_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_247_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_248_clock; // @[mac.scala 29:63]
  wire  PECross_248_reset; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_248_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_248_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_248_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_248_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_248_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_248_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_248_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_248_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_249_clock; // @[mac.scala 29:63]
  wire  PECross_249_reset; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_249_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_249_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_249_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_249_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_249_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_249_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_249_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_249_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_250_clock; // @[mac.scala 29:63]
  wire  PECross_250_reset; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_250_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_250_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_250_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_250_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_250_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_250_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_250_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_250_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_251_clock; // @[mac.scala 29:63]
  wire  PECross_251_reset; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_251_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_251_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_251_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_251_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_251_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_251_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_251_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_251_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_252_clock; // @[mac.scala 29:63]
  wire  PECross_252_reset; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_252_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_252_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_252_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_252_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_252_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_252_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_252_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_252_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_253_clock; // @[mac.scala 29:63]
  wire  PECross_253_reset; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_253_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_253_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_253_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_253_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_253_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_253_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_253_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_253_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_254_clock; // @[mac.scala 29:63]
  wire  PECross_254_reset; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_254_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_254_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_254_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_254_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_254_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_254_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_254_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_254_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_255_clock; // @[mac.scala 29:63]
  wire  PECross_255_reset; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_sumIn_ready; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_sumIn_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_255_multiply_io_input_io_sumIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_sumIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_sumOut_ready; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_sumOut_valid; // @[mac.scala 29:63]
  wire [19:0] PECross_255_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 29:63]
  wire [1:0] PECross_255_multiply_io_input_io_statSel; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiEn; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actEn; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actIn_ready; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_255_multiply_io_input_io_actIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiIn_ready; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiIn_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_255_multiply_io_input_io_weiIn_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiIn_bits_last; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actOut_ready; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_255_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_actOut_bits_last; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiOut_ready; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiOut_valid; // @[mac.scala 29:63]
  wire [7:0] PECross_255_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 29:63]
  wire  PECross_255_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 29:63]
  PECross PECross ( // @[mac.scala 29:63]
    .clock(PECross_clock),
    .reset(PECross_reset),
    .multiply_io_input_io_sumIn_ready(PECross_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_1 ( // @[mac.scala 29:63]
    .clock(PECross_1_clock),
    .reset(PECross_1_reset),
    .multiply_io_input_io_sumIn_ready(PECross_1_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_1_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_1_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_1_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_1_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_1_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_1_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_1_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_1_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_1_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_1_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_1_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_1_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_1_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_1_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_1_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_1_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_1_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_1_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_1_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_1_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_1_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_1_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_1_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_1_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_1_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_1_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_2 ( // @[mac.scala 29:63]
    .clock(PECross_2_clock),
    .reset(PECross_2_reset),
    .multiply_io_input_io_sumIn_ready(PECross_2_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_2_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_2_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_2_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_2_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_2_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_2_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_2_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_2_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_2_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_2_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_2_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_2_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_2_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_2_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_2_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_2_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_2_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_2_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_2_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_2_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_2_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_2_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_2_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_2_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_2_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_2_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_3 ( // @[mac.scala 29:63]
    .clock(PECross_3_clock),
    .reset(PECross_3_reset),
    .multiply_io_input_io_sumIn_ready(PECross_3_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_3_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_3_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_3_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_3_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_3_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_3_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_3_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_3_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_3_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_3_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_3_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_3_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_3_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_3_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_3_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_3_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_3_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_3_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_3_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_3_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_3_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_3_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_3_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_3_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_3_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_3_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_4 ( // @[mac.scala 29:63]
    .clock(PECross_4_clock),
    .reset(PECross_4_reset),
    .multiply_io_input_io_sumIn_ready(PECross_4_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_4_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_4_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_4_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_4_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_4_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_4_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_4_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_4_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_4_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_4_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_4_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_4_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_4_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_4_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_4_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_4_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_4_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_4_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_4_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_4_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_4_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_4_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_4_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_4_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_4_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_4_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_5 ( // @[mac.scala 29:63]
    .clock(PECross_5_clock),
    .reset(PECross_5_reset),
    .multiply_io_input_io_sumIn_ready(PECross_5_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_5_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_5_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_5_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_5_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_5_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_5_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_5_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_5_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_5_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_5_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_5_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_5_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_5_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_5_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_5_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_5_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_5_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_5_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_5_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_5_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_5_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_5_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_5_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_5_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_5_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_5_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_6 ( // @[mac.scala 29:63]
    .clock(PECross_6_clock),
    .reset(PECross_6_reset),
    .multiply_io_input_io_sumIn_ready(PECross_6_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_6_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_6_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_6_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_6_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_6_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_6_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_6_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_6_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_6_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_6_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_6_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_6_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_6_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_6_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_6_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_6_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_6_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_6_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_6_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_6_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_6_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_6_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_6_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_6_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_6_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_6_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_7 ( // @[mac.scala 29:63]
    .clock(PECross_7_clock),
    .reset(PECross_7_reset),
    .multiply_io_input_io_sumIn_ready(PECross_7_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_7_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_7_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_7_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_7_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_7_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_7_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_7_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_7_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_7_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_7_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_7_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_7_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_7_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_7_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_7_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_7_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_7_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_7_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_7_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_7_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_7_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_7_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_7_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_7_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_7_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_7_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_8 ( // @[mac.scala 29:63]
    .clock(PECross_8_clock),
    .reset(PECross_8_reset),
    .multiply_io_input_io_sumIn_ready(PECross_8_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_8_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_8_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_8_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_8_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_8_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_8_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_8_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_8_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_8_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_8_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_8_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_8_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_8_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_8_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_8_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_8_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_8_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_8_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_8_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_8_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_8_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_8_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_8_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_8_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_8_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_8_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_9 ( // @[mac.scala 29:63]
    .clock(PECross_9_clock),
    .reset(PECross_9_reset),
    .multiply_io_input_io_sumIn_ready(PECross_9_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_9_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_9_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_9_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_9_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_9_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_9_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_9_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_9_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_9_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_9_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_9_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_9_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_9_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_9_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_9_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_9_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_9_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_9_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_9_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_9_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_9_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_9_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_9_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_9_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_9_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_9_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_10 ( // @[mac.scala 29:63]
    .clock(PECross_10_clock),
    .reset(PECross_10_reset),
    .multiply_io_input_io_sumIn_ready(PECross_10_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_10_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_10_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_10_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_10_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_10_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_10_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_10_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_10_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_10_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_10_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_10_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_10_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_10_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_10_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_10_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_10_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_10_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_10_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_10_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_10_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_10_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_10_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_10_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_10_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_10_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_10_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_11 ( // @[mac.scala 29:63]
    .clock(PECross_11_clock),
    .reset(PECross_11_reset),
    .multiply_io_input_io_sumIn_ready(PECross_11_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_11_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_11_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_11_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_11_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_11_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_11_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_11_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_11_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_11_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_11_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_11_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_11_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_11_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_11_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_11_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_11_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_11_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_11_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_11_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_11_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_11_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_11_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_11_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_11_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_11_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_11_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_12 ( // @[mac.scala 29:63]
    .clock(PECross_12_clock),
    .reset(PECross_12_reset),
    .multiply_io_input_io_sumIn_ready(PECross_12_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_12_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_12_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_12_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_12_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_12_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_12_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_12_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_12_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_12_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_12_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_12_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_12_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_12_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_12_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_12_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_12_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_12_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_12_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_12_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_12_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_12_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_12_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_12_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_12_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_12_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_12_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_13 ( // @[mac.scala 29:63]
    .clock(PECross_13_clock),
    .reset(PECross_13_reset),
    .multiply_io_input_io_sumIn_ready(PECross_13_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_13_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_13_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_13_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_13_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_13_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_13_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_13_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_13_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_13_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_13_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_13_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_13_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_13_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_13_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_13_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_13_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_13_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_13_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_13_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_13_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_13_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_13_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_13_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_13_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_13_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_13_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_14 ( // @[mac.scala 29:63]
    .clock(PECross_14_clock),
    .reset(PECross_14_reset),
    .multiply_io_input_io_sumIn_ready(PECross_14_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_14_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_14_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_14_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_14_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_14_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_14_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_14_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_14_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_14_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_14_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_14_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_14_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_14_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_14_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_14_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_14_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_14_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_14_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_14_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_14_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_14_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_14_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_14_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_14_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_14_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_14_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_15 ( // @[mac.scala 29:63]
    .clock(PECross_15_clock),
    .reset(PECross_15_reset),
    .multiply_io_input_io_sumIn_ready(PECross_15_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_15_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_15_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_15_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_15_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_15_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_15_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_15_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_15_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_15_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_15_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_15_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_15_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_15_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_15_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_15_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_15_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_15_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_15_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_15_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_15_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_15_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_15_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_15_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_15_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_15_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_15_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_16 ( // @[mac.scala 29:63]
    .clock(PECross_16_clock),
    .reset(PECross_16_reset),
    .multiply_io_input_io_sumIn_ready(PECross_16_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_16_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_16_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_16_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_16_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_16_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_16_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_16_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_16_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_16_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_16_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_16_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_16_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_16_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_16_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_16_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_16_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_16_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_16_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_16_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_16_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_16_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_16_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_16_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_16_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_16_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_16_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_17 ( // @[mac.scala 29:63]
    .clock(PECross_17_clock),
    .reset(PECross_17_reset),
    .multiply_io_input_io_sumIn_ready(PECross_17_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_17_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_17_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_17_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_17_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_17_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_17_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_17_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_17_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_17_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_17_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_17_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_17_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_17_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_17_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_17_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_17_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_17_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_17_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_17_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_17_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_17_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_17_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_17_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_17_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_17_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_17_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_18 ( // @[mac.scala 29:63]
    .clock(PECross_18_clock),
    .reset(PECross_18_reset),
    .multiply_io_input_io_sumIn_ready(PECross_18_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_18_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_18_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_18_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_18_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_18_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_18_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_18_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_18_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_18_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_18_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_18_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_18_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_18_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_18_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_18_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_18_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_18_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_18_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_18_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_18_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_18_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_18_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_18_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_18_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_18_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_18_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_19 ( // @[mac.scala 29:63]
    .clock(PECross_19_clock),
    .reset(PECross_19_reset),
    .multiply_io_input_io_sumIn_ready(PECross_19_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_19_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_19_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_19_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_19_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_19_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_19_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_19_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_19_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_19_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_19_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_19_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_19_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_19_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_19_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_19_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_19_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_19_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_19_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_19_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_19_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_19_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_19_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_19_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_19_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_19_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_19_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_20 ( // @[mac.scala 29:63]
    .clock(PECross_20_clock),
    .reset(PECross_20_reset),
    .multiply_io_input_io_sumIn_ready(PECross_20_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_20_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_20_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_20_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_20_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_20_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_20_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_20_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_20_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_20_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_20_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_20_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_20_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_20_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_20_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_20_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_20_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_20_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_20_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_20_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_20_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_20_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_20_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_20_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_20_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_20_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_20_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_21 ( // @[mac.scala 29:63]
    .clock(PECross_21_clock),
    .reset(PECross_21_reset),
    .multiply_io_input_io_sumIn_ready(PECross_21_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_21_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_21_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_21_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_21_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_21_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_21_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_21_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_21_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_21_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_21_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_21_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_21_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_21_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_21_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_21_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_21_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_21_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_21_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_21_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_21_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_21_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_21_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_21_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_21_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_21_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_21_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_22 ( // @[mac.scala 29:63]
    .clock(PECross_22_clock),
    .reset(PECross_22_reset),
    .multiply_io_input_io_sumIn_ready(PECross_22_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_22_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_22_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_22_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_22_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_22_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_22_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_22_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_22_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_22_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_22_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_22_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_22_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_22_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_22_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_22_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_22_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_22_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_22_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_22_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_22_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_22_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_22_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_22_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_22_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_22_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_22_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_23 ( // @[mac.scala 29:63]
    .clock(PECross_23_clock),
    .reset(PECross_23_reset),
    .multiply_io_input_io_sumIn_ready(PECross_23_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_23_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_23_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_23_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_23_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_23_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_23_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_23_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_23_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_23_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_23_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_23_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_23_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_23_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_23_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_23_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_23_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_23_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_23_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_23_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_23_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_23_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_23_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_23_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_23_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_23_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_23_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_24 ( // @[mac.scala 29:63]
    .clock(PECross_24_clock),
    .reset(PECross_24_reset),
    .multiply_io_input_io_sumIn_ready(PECross_24_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_24_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_24_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_24_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_24_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_24_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_24_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_24_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_24_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_24_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_24_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_24_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_24_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_24_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_24_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_24_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_24_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_24_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_24_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_24_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_24_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_24_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_24_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_24_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_24_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_24_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_24_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_25 ( // @[mac.scala 29:63]
    .clock(PECross_25_clock),
    .reset(PECross_25_reset),
    .multiply_io_input_io_sumIn_ready(PECross_25_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_25_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_25_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_25_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_25_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_25_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_25_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_25_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_25_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_25_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_25_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_25_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_25_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_25_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_25_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_25_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_25_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_25_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_25_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_25_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_25_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_25_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_25_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_25_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_25_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_25_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_25_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_26 ( // @[mac.scala 29:63]
    .clock(PECross_26_clock),
    .reset(PECross_26_reset),
    .multiply_io_input_io_sumIn_ready(PECross_26_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_26_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_26_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_26_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_26_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_26_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_26_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_26_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_26_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_26_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_26_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_26_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_26_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_26_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_26_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_26_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_26_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_26_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_26_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_26_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_26_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_26_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_26_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_26_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_26_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_26_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_26_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_27 ( // @[mac.scala 29:63]
    .clock(PECross_27_clock),
    .reset(PECross_27_reset),
    .multiply_io_input_io_sumIn_ready(PECross_27_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_27_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_27_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_27_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_27_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_27_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_27_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_27_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_27_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_27_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_27_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_27_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_27_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_27_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_27_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_27_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_27_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_27_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_27_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_27_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_27_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_27_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_27_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_27_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_27_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_27_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_27_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_28 ( // @[mac.scala 29:63]
    .clock(PECross_28_clock),
    .reset(PECross_28_reset),
    .multiply_io_input_io_sumIn_ready(PECross_28_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_28_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_28_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_28_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_28_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_28_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_28_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_28_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_28_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_28_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_28_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_28_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_28_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_28_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_28_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_28_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_28_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_28_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_28_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_28_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_28_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_28_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_28_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_28_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_28_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_28_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_28_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_29 ( // @[mac.scala 29:63]
    .clock(PECross_29_clock),
    .reset(PECross_29_reset),
    .multiply_io_input_io_sumIn_ready(PECross_29_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_29_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_29_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_29_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_29_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_29_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_29_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_29_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_29_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_29_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_29_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_29_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_29_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_29_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_29_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_29_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_29_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_29_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_29_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_29_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_29_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_29_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_29_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_29_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_29_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_29_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_29_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_30 ( // @[mac.scala 29:63]
    .clock(PECross_30_clock),
    .reset(PECross_30_reset),
    .multiply_io_input_io_sumIn_ready(PECross_30_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_30_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_30_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_30_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_30_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_30_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_30_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_30_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_30_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_30_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_30_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_30_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_30_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_30_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_30_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_30_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_30_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_30_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_30_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_30_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_30_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_30_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_30_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_30_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_30_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_30_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_30_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_31 ( // @[mac.scala 29:63]
    .clock(PECross_31_clock),
    .reset(PECross_31_reset),
    .multiply_io_input_io_sumIn_ready(PECross_31_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_31_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_31_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_31_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_31_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_31_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_31_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_31_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_31_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_31_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_31_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_31_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_31_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_31_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_31_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_31_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_31_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_31_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_31_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_31_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_31_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_31_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_31_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_31_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_31_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_31_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_31_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_32 ( // @[mac.scala 29:63]
    .clock(PECross_32_clock),
    .reset(PECross_32_reset),
    .multiply_io_input_io_sumIn_ready(PECross_32_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_32_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_32_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_32_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_32_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_32_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_32_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_32_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_32_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_32_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_32_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_32_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_32_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_32_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_32_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_32_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_32_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_32_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_32_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_32_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_32_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_32_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_32_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_32_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_32_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_32_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_32_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_33 ( // @[mac.scala 29:63]
    .clock(PECross_33_clock),
    .reset(PECross_33_reset),
    .multiply_io_input_io_sumIn_ready(PECross_33_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_33_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_33_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_33_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_33_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_33_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_33_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_33_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_33_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_33_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_33_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_33_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_33_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_33_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_33_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_33_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_33_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_33_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_33_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_33_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_33_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_33_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_33_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_33_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_33_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_33_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_33_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_34 ( // @[mac.scala 29:63]
    .clock(PECross_34_clock),
    .reset(PECross_34_reset),
    .multiply_io_input_io_sumIn_ready(PECross_34_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_34_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_34_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_34_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_34_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_34_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_34_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_34_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_34_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_34_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_34_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_34_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_34_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_34_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_34_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_34_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_34_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_34_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_34_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_34_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_34_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_34_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_34_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_34_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_34_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_34_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_34_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_35 ( // @[mac.scala 29:63]
    .clock(PECross_35_clock),
    .reset(PECross_35_reset),
    .multiply_io_input_io_sumIn_ready(PECross_35_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_35_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_35_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_35_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_35_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_35_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_35_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_35_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_35_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_35_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_35_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_35_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_35_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_35_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_35_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_35_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_35_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_35_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_35_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_35_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_35_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_35_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_35_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_35_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_35_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_35_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_35_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_36 ( // @[mac.scala 29:63]
    .clock(PECross_36_clock),
    .reset(PECross_36_reset),
    .multiply_io_input_io_sumIn_ready(PECross_36_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_36_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_36_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_36_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_36_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_36_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_36_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_36_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_36_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_36_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_36_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_36_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_36_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_36_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_36_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_36_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_36_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_36_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_36_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_36_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_36_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_36_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_36_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_36_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_36_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_36_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_36_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_37 ( // @[mac.scala 29:63]
    .clock(PECross_37_clock),
    .reset(PECross_37_reset),
    .multiply_io_input_io_sumIn_ready(PECross_37_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_37_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_37_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_37_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_37_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_37_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_37_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_37_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_37_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_37_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_37_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_37_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_37_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_37_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_37_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_37_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_37_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_37_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_37_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_37_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_37_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_37_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_37_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_37_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_37_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_37_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_37_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_38 ( // @[mac.scala 29:63]
    .clock(PECross_38_clock),
    .reset(PECross_38_reset),
    .multiply_io_input_io_sumIn_ready(PECross_38_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_38_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_38_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_38_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_38_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_38_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_38_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_38_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_38_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_38_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_38_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_38_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_38_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_38_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_38_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_38_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_38_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_38_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_38_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_38_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_38_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_38_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_38_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_38_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_38_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_38_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_38_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_39 ( // @[mac.scala 29:63]
    .clock(PECross_39_clock),
    .reset(PECross_39_reset),
    .multiply_io_input_io_sumIn_ready(PECross_39_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_39_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_39_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_39_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_39_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_39_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_39_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_39_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_39_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_39_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_39_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_39_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_39_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_39_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_39_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_39_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_39_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_39_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_39_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_39_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_39_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_39_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_39_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_39_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_39_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_39_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_39_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_40 ( // @[mac.scala 29:63]
    .clock(PECross_40_clock),
    .reset(PECross_40_reset),
    .multiply_io_input_io_sumIn_ready(PECross_40_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_40_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_40_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_40_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_40_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_40_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_40_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_40_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_40_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_40_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_40_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_40_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_40_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_40_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_40_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_40_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_40_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_40_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_40_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_40_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_40_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_40_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_40_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_40_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_40_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_40_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_40_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_41 ( // @[mac.scala 29:63]
    .clock(PECross_41_clock),
    .reset(PECross_41_reset),
    .multiply_io_input_io_sumIn_ready(PECross_41_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_41_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_41_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_41_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_41_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_41_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_41_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_41_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_41_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_41_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_41_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_41_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_41_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_41_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_41_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_41_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_41_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_41_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_41_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_41_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_41_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_41_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_41_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_41_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_41_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_41_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_41_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_42 ( // @[mac.scala 29:63]
    .clock(PECross_42_clock),
    .reset(PECross_42_reset),
    .multiply_io_input_io_sumIn_ready(PECross_42_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_42_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_42_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_42_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_42_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_42_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_42_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_42_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_42_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_42_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_42_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_42_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_42_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_42_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_42_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_42_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_42_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_42_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_42_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_42_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_42_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_42_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_42_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_42_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_42_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_42_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_42_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_43 ( // @[mac.scala 29:63]
    .clock(PECross_43_clock),
    .reset(PECross_43_reset),
    .multiply_io_input_io_sumIn_ready(PECross_43_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_43_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_43_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_43_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_43_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_43_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_43_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_43_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_43_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_43_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_43_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_43_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_43_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_43_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_43_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_43_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_43_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_43_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_43_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_43_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_43_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_43_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_43_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_43_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_43_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_43_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_43_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_44 ( // @[mac.scala 29:63]
    .clock(PECross_44_clock),
    .reset(PECross_44_reset),
    .multiply_io_input_io_sumIn_ready(PECross_44_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_44_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_44_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_44_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_44_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_44_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_44_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_44_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_44_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_44_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_44_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_44_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_44_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_44_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_44_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_44_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_44_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_44_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_44_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_44_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_44_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_44_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_44_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_44_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_44_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_44_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_44_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_45 ( // @[mac.scala 29:63]
    .clock(PECross_45_clock),
    .reset(PECross_45_reset),
    .multiply_io_input_io_sumIn_ready(PECross_45_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_45_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_45_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_45_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_45_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_45_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_45_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_45_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_45_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_45_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_45_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_45_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_45_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_45_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_45_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_45_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_45_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_45_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_45_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_45_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_45_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_45_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_45_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_45_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_45_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_45_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_45_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_46 ( // @[mac.scala 29:63]
    .clock(PECross_46_clock),
    .reset(PECross_46_reset),
    .multiply_io_input_io_sumIn_ready(PECross_46_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_46_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_46_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_46_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_46_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_46_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_46_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_46_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_46_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_46_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_46_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_46_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_46_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_46_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_46_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_46_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_46_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_46_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_46_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_46_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_46_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_46_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_46_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_46_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_46_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_46_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_46_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_47 ( // @[mac.scala 29:63]
    .clock(PECross_47_clock),
    .reset(PECross_47_reset),
    .multiply_io_input_io_sumIn_ready(PECross_47_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_47_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_47_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_47_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_47_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_47_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_47_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_47_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_47_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_47_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_47_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_47_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_47_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_47_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_47_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_47_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_47_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_47_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_47_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_47_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_47_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_47_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_47_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_47_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_47_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_47_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_47_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_48 ( // @[mac.scala 29:63]
    .clock(PECross_48_clock),
    .reset(PECross_48_reset),
    .multiply_io_input_io_sumIn_ready(PECross_48_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_48_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_48_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_48_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_48_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_48_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_48_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_48_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_48_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_48_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_48_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_48_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_48_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_48_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_48_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_48_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_48_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_48_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_48_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_48_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_48_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_48_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_48_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_48_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_48_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_48_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_48_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_49 ( // @[mac.scala 29:63]
    .clock(PECross_49_clock),
    .reset(PECross_49_reset),
    .multiply_io_input_io_sumIn_ready(PECross_49_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_49_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_49_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_49_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_49_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_49_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_49_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_49_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_49_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_49_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_49_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_49_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_49_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_49_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_49_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_49_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_49_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_49_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_49_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_49_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_49_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_49_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_49_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_49_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_49_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_49_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_49_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_50 ( // @[mac.scala 29:63]
    .clock(PECross_50_clock),
    .reset(PECross_50_reset),
    .multiply_io_input_io_sumIn_ready(PECross_50_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_50_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_50_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_50_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_50_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_50_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_50_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_50_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_50_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_50_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_50_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_50_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_50_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_50_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_50_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_50_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_50_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_50_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_50_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_50_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_50_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_50_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_50_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_50_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_50_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_50_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_50_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_51 ( // @[mac.scala 29:63]
    .clock(PECross_51_clock),
    .reset(PECross_51_reset),
    .multiply_io_input_io_sumIn_ready(PECross_51_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_51_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_51_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_51_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_51_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_51_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_51_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_51_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_51_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_51_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_51_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_51_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_51_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_51_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_51_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_51_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_51_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_51_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_51_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_51_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_51_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_51_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_51_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_51_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_51_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_51_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_51_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_52 ( // @[mac.scala 29:63]
    .clock(PECross_52_clock),
    .reset(PECross_52_reset),
    .multiply_io_input_io_sumIn_ready(PECross_52_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_52_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_52_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_52_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_52_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_52_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_52_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_52_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_52_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_52_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_52_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_52_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_52_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_52_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_52_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_52_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_52_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_52_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_52_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_52_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_52_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_52_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_52_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_52_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_52_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_52_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_52_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_53 ( // @[mac.scala 29:63]
    .clock(PECross_53_clock),
    .reset(PECross_53_reset),
    .multiply_io_input_io_sumIn_ready(PECross_53_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_53_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_53_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_53_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_53_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_53_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_53_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_53_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_53_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_53_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_53_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_53_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_53_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_53_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_53_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_53_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_53_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_53_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_53_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_53_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_53_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_53_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_53_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_53_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_53_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_53_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_53_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_54 ( // @[mac.scala 29:63]
    .clock(PECross_54_clock),
    .reset(PECross_54_reset),
    .multiply_io_input_io_sumIn_ready(PECross_54_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_54_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_54_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_54_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_54_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_54_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_54_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_54_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_54_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_54_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_54_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_54_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_54_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_54_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_54_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_54_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_54_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_54_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_54_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_54_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_54_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_54_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_54_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_54_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_54_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_54_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_54_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_55 ( // @[mac.scala 29:63]
    .clock(PECross_55_clock),
    .reset(PECross_55_reset),
    .multiply_io_input_io_sumIn_ready(PECross_55_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_55_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_55_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_55_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_55_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_55_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_55_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_55_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_55_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_55_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_55_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_55_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_55_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_55_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_55_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_55_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_55_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_55_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_55_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_55_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_55_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_55_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_55_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_55_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_55_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_55_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_55_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_56 ( // @[mac.scala 29:63]
    .clock(PECross_56_clock),
    .reset(PECross_56_reset),
    .multiply_io_input_io_sumIn_ready(PECross_56_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_56_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_56_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_56_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_56_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_56_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_56_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_56_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_56_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_56_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_56_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_56_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_56_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_56_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_56_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_56_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_56_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_56_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_56_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_56_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_56_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_56_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_56_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_56_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_56_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_56_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_56_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_57 ( // @[mac.scala 29:63]
    .clock(PECross_57_clock),
    .reset(PECross_57_reset),
    .multiply_io_input_io_sumIn_ready(PECross_57_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_57_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_57_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_57_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_57_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_57_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_57_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_57_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_57_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_57_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_57_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_57_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_57_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_57_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_57_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_57_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_57_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_57_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_57_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_57_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_57_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_57_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_57_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_57_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_57_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_57_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_57_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_58 ( // @[mac.scala 29:63]
    .clock(PECross_58_clock),
    .reset(PECross_58_reset),
    .multiply_io_input_io_sumIn_ready(PECross_58_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_58_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_58_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_58_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_58_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_58_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_58_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_58_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_58_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_58_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_58_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_58_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_58_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_58_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_58_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_58_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_58_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_58_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_58_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_58_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_58_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_58_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_58_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_58_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_58_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_58_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_58_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_59 ( // @[mac.scala 29:63]
    .clock(PECross_59_clock),
    .reset(PECross_59_reset),
    .multiply_io_input_io_sumIn_ready(PECross_59_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_59_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_59_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_59_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_59_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_59_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_59_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_59_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_59_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_59_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_59_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_59_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_59_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_59_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_59_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_59_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_59_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_59_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_59_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_59_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_59_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_59_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_59_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_59_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_59_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_59_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_59_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_60 ( // @[mac.scala 29:63]
    .clock(PECross_60_clock),
    .reset(PECross_60_reset),
    .multiply_io_input_io_sumIn_ready(PECross_60_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_60_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_60_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_60_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_60_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_60_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_60_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_60_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_60_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_60_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_60_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_60_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_60_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_60_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_60_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_60_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_60_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_60_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_60_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_60_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_60_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_60_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_60_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_60_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_60_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_60_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_60_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_61 ( // @[mac.scala 29:63]
    .clock(PECross_61_clock),
    .reset(PECross_61_reset),
    .multiply_io_input_io_sumIn_ready(PECross_61_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_61_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_61_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_61_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_61_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_61_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_61_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_61_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_61_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_61_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_61_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_61_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_61_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_61_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_61_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_61_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_61_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_61_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_61_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_61_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_61_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_61_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_61_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_61_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_61_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_61_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_61_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_62 ( // @[mac.scala 29:63]
    .clock(PECross_62_clock),
    .reset(PECross_62_reset),
    .multiply_io_input_io_sumIn_ready(PECross_62_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_62_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_62_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_62_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_62_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_62_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_62_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_62_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_62_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_62_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_62_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_62_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_62_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_62_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_62_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_62_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_62_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_62_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_62_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_62_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_62_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_62_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_62_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_62_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_62_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_62_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_62_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_63 ( // @[mac.scala 29:63]
    .clock(PECross_63_clock),
    .reset(PECross_63_reset),
    .multiply_io_input_io_sumIn_ready(PECross_63_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_63_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_63_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_63_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_63_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_63_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_63_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_63_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_63_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_63_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_63_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_63_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_63_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_63_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_63_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_63_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_63_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_63_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_63_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_63_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_63_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_63_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_63_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_63_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_63_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_63_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_63_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_64 ( // @[mac.scala 29:63]
    .clock(PECross_64_clock),
    .reset(PECross_64_reset),
    .multiply_io_input_io_sumIn_ready(PECross_64_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_64_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_64_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_64_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_64_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_64_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_64_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_64_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_64_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_64_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_64_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_64_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_64_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_64_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_64_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_64_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_64_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_64_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_64_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_64_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_64_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_64_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_64_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_64_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_64_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_64_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_64_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_65 ( // @[mac.scala 29:63]
    .clock(PECross_65_clock),
    .reset(PECross_65_reset),
    .multiply_io_input_io_sumIn_ready(PECross_65_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_65_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_65_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_65_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_65_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_65_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_65_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_65_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_65_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_65_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_65_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_65_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_65_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_65_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_65_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_65_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_65_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_65_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_65_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_65_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_65_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_65_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_65_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_65_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_65_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_65_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_65_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_66 ( // @[mac.scala 29:63]
    .clock(PECross_66_clock),
    .reset(PECross_66_reset),
    .multiply_io_input_io_sumIn_ready(PECross_66_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_66_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_66_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_66_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_66_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_66_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_66_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_66_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_66_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_66_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_66_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_66_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_66_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_66_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_66_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_66_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_66_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_66_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_66_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_66_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_66_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_66_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_66_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_66_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_66_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_66_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_66_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_67 ( // @[mac.scala 29:63]
    .clock(PECross_67_clock),
    .reset(PECross_67_reset),
    .multiply_io_input_io_sumIn_ready(PECross_67_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_67_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_67_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_67_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_67_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_67_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_67_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_67_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_67_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_67_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_67_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_67_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_67_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_67_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_67_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_67_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_67_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_67_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_67_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_67_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_67_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_67_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_67_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_67_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_67_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_67_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_67_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_68 ( // @[mac.scala 29:63]
    .clock(PECross_68_clock),
    .reset(PECross_68_reset),
    .multiply_io_input_io_sumIn_ready(PECross_68_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_68_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_68_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_68_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_68_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_68_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_68_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_68_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_68_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_68_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_68_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_68_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_68_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_68_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_68_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_68_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_68_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_68_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_68_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_68_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_68_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_68_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_68_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_68_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_68_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_68_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_68_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_69 ( // @[mac.scala 29:63]
    .clock(PECross_69_clock),
    .reset(PECross_69_reset),
    .multiply_io_input_io_sumIn_ready(PECross_69_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_69_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_69_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_69_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_69_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_69_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_69_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_69_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_69_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_69_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_69_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_69_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_69_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_69_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_69_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_69_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_69_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_69_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_69_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_69_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_69_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_69_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_69_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_69_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_69_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_69_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_69_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_70 ( // @[mac.scala 29:63]
    .clock(PECross_70_clock),
    .reset(PECross_70_reset),
    .multiply_io_input_io_sumIn_ready(PECross_70_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_70_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_70_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_70_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_70_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_70_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_70_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_70_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_70_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_70_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_70_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_70_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_70_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_70_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_70_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_70_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_70_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_70_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_70_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_70_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_70_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_70_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_70_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_70_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_70_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_70_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_70_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_71 ( // @[mac.scala 29:63]
    .clock(PECross_71_clock),
    .reset(PECross_71_reset),
    .multiply_io_input_io_sumIn_ready(PECross_71_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_71_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_71_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_71_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_71_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_71_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_71_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_71_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_71_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_71_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_71_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_71_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_71_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_71_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_71_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_71_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_71_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_71_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_71_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_71_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_71_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_71_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_71_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_71_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_71_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_71_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_71_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_72 ( // @[mac.scala 29:63]
    .clock(PECross_72_clock),
    .reset(PECross_72_reset),
    .multiply_io_input_io_sumIn_ready(PECross_72_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_72_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_72_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_72_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_72_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_72_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_72_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_72_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_72_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_72_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_72_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_72_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_72_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_72_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_72_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_72_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_72_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_72_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_72_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_72_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_72_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_72_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_72_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_72_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_72_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_72_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_72_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_73 ( // @[mac.scala 29:63]
    .clock(PECross_73_clock),
    .reset(PECross_73_reset),
    .multiply_io_input_io_sumIn_ready(PECross_73_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_73_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_73_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_73_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_73_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_73_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_73_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_73_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_73_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_73_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_73_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_73_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_73_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_73_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_73_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_73_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_73_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_73_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_73_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_73_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_73_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_73_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_73_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_73_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_73_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_73_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_73_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_74 ( // @[mac.scala 29:63]
    .clock(PECross_74_clock),
    .reset(PECross_74_reset),
    .multiply_io_input_io_sumIn_ready(PECross_74_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_74_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_74_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_74_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_74_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_74_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_74_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_74_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_74_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_74_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_74_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_74_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_74_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_74_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_74_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_74_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_74_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_74_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_74_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_74_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_74_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_74_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_74_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_74_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_74_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_74_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_74_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_75 ( // @[mac.scala 29:63]
    .clock(PECross_75_clock),
    .reset(PECross_75_reset),
    .multiply_io_input_io_sumIn_ready(PECross_75_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_75_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_75_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_75_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_75_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_75_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_75_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_75_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_75_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_75_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_75_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_75_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_75_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_75_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_75_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_75_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_75_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_75_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_75_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_75_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_75_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_75_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_75_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_75_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_75_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_75_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_75_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_76 ( // @[mac.scala 29:63]
    .clock(PECross_76_clock),
    .reset(PECross_76_reset),
    .multiply_io_input_io_sumIn_ready(PECross_76_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_76_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_76_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_76_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_76_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_76_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_76_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_76_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_76_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_76_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_76_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_76_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_76_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_76_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_76_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_76_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_76_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_76_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_76_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_76_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_76_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_76_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_76_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_76_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_76_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_76_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_76_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_77 ( // @[mac.scala 29:63]
    .clock(PECross_77_clock),
    .reset(PECross_77_reset),
    .multiply_io_input_io_sumIn_ready(PECross_77_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_77_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_77_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_77_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_77_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_77_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_77_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_77_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_77_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_77_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_77_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_77_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_77_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_77_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_77_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_77_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_77_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_77_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_77_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_77_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_77_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_77_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_77_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_77_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_77_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_77_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_77_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_78 ( // @[mac.scala 29:63]
    .clock(PECross_78_clock),
    .reset(PECross_78_reset),
    .multiply_io_input_io_sumIn_ready(PECross_78_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_78_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_78_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_78_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_78_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_78_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_78_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_78_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_78_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_78_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_78_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_78_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_78_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_78_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_78_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_78_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_78_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_78_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_78_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_78_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_78_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_78_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_78_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_78_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_78_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_78_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_78_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_79 ( // @[mac.scala 29:63]
    .clock(PECross_79_clock),
    .reset(PECross_79_reset),
    .multiply_io_input_io_sumIn_ready(PECross_79_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_79_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_79_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_79_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_79_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_79_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_79_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_79_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_79_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_79_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_79_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_79_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_79_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_79_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_79_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_79_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_79_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_79_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_79_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_79_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_79_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_79_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_79_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_79_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_79_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_79_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_79_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_80 ( // @[mac.scala 29:63]
    .clock(PECross_80_clock),
    .reset(PECross_80_reset),
    .multiply_io_input_io_sumIn_ready(PECross_80_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_80_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_80_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_80_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_80_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_80_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_80_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_80_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_80_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_80_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_80_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_80_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_80_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_80_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_80_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_80_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_80_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_80_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_80_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_80_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_80_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_80_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_80_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_80_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_80_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_80_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_80_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_81 ( // @[mac.scala 29:63]
    .clock(PECross_81_clock),
    .reset(PECross_81_reset),
    .multiply_io_input_io_sumIn_ready(PECross_81_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_81_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_81_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_81_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_81_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_81_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_81_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_81_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_81_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_81_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_81_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_81_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_81_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_81_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_81_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_81_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_81_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_81_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_81_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_81_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_81_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_81_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_81_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_81_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_81_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_81_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_81_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_82 ( // @[mac.scala 29:63]
    .clock(PECross_82_clock),
    .reset(PECross_82_reset),
    .multiply_io_input_io_sumIn_ready(PECross_82_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_82_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_82_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_82_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_82_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_82_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_82_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_82_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_82_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_82_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_82_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_82_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_82_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_82_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_82_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_82_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_82_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_82_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_82_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_82_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_82_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_82_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_82_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_82_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_82_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_82_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_82_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_83 ( // @[mac.scala 29:63]
    .clock(PECross_83_clock),
    .reset(PECross_83_reset),
    .multiply_io_input_io_sumIn_ready(PECross_83_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_83_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_83_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_83_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_83_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_83_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_83_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_83_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_83_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_83_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_83_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_83_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_83_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_83_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_83_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_83_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_83_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_83_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_83_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_83_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_83_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_83_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_83_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_83_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_83_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_83_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_83_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_84 ( // @[mac.scala 29:63]
    .clock(PECross_84_clock),
    .reset(PECross_84_reset),
    .multiply_io_input_io_sumIn_ready(PECross_84_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_84_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_84_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_84_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_84_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_84_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_84_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_84_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_84_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_84_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_84_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_84_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_84_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_84_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_84_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_84_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_84_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_84_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_84_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_84_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_84_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_84_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_84_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_84_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_84_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_84_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_84_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_85 ( // @[mac.scala 29:63]
    .clock(PECross_85_clock),
    .reset(PECross_85_reset),
    .multiply_io_input_io_sumIn_ready(PECross_85_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_85_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_85_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_85_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_85_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_85_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_85_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_85_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_85_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_85_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_85_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_85_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_85_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_85_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_85_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_85_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_85_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_85_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_85_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_85_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_85_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_85_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_85_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_85_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_85_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_85_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_85_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_86 ( // @[mac.scala 29:63]
    .clock(PECross_86_clock),
    .reset(PECross_86_reset),
    .multiply_io_input_io_sumIn_ready(PECross_86_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_86_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_86_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_86_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_86_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_86_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_86_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_86_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_86_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_86_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_86_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_86_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_86_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_86_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_86_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_86_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_86_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_86_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_86_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_86_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_86_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_86_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_86_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_86_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_86_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_86_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_86_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_87 ( // @[mac.scala 29:63]
    .clock(PECross_87_clock),
    .reset(PECross_87_reset),
    .multiply_io_input_io_sumIn_ready(PECross_87_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_87_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_87_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_87_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_87_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_87_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_87_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_87_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_87_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_87_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_87_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_87_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_87_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_87_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_87_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_87_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_87_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_87_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_87_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_87_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_87_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_87_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_87_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_87_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_87_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_87_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_87_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_88 ( // @[mac.scala 29:63]
    .clock(PECross_88_clock),
    .reset(PECross_88_reset),
    .multiply_io_input_io_sumIn_ready(PECross_88_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_88_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_88_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_88_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_88_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_88_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_88_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_88_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_88_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_88_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_88_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_88_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_88_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_88_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_88_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_88_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_88_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_88_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_88_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_88_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_88_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_88_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_88_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_88_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_88_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_88_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_88_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_89 ( // @[mac.scala 29:63]
    .clock(PECross_89_clock),
    .reset(PECross_89_reset),
    .multiply_io_input_io_sumIn_ready(PECross_89_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_89_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_89_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_89_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_89_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_89_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_89_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_89_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_89_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_89_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_89_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_89_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_89_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_89_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_89_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_89_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_89_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_89_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_89_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_89_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_89_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_89_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_89_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_89_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_89_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_89_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_89_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_90 ( // @[mac.scala 29:63]
    .clock(PECross_90_clock),
    .reset(PECross_90_reset),
    .multiply_io_input_io_sumIn_ready(PECross_90_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_90_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_90_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_90_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_90_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_90_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_90_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_90_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_90_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_90_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_90_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_90_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_90_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_90_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_90_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_90_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_90_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_90_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_90_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_90_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_90_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_90_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_90_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_90_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_90_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_90_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_90_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_91 ( // @[mac.scala 29:63]
    .clock(PECross_91_clock),
    .reset(PECross_91_reset),
    .multiply_io_input_io_sumIn_ready(PECross_91_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_91_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_91_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_91_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_91_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_91_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_91_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_91_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_91_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_91_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_91_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_91_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_91_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_91_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_91_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_91_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_91_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_91_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_91_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_91_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_91_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_91_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_91_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_91_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_91_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_91_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_91_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_92 ( // @[mac.scala 29:63]
    .clock(PECross_92_clock),
    .reset(PECross_92_reset),
    .multiply_io_input_io_sumIn_ready(PECross_92_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_92_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_92_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_92_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_92_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_92_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_92_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_92_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_92_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_92_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_92_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_92_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_92_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_92_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_92_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_92_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_92_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_92_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_92_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_92_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_92_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_92_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_92_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_92_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_92_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_92_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_92_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_93 ( // @[mac.scala 29:63]
    .clock(PECross_93_clock),
    .reset(PECross_93_reset),
    .multiply_io_input_io_sumIn_ready(PECross_93_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_93_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_93_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_93_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_93_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_93_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_93_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_93_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_93_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_93_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_93_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_93_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_93_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_93_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_93_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_93_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_93_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_93_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_93_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_93_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_93_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_93_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_93_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_93_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_93_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_93_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_93_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_94 ( // @[mac.scala 29:63]
    .clock(PECross_94_clock),
    .reset(PECross_94_reset),
    .multiply_io_input_io_sumIn_ready(PECross_94_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_94_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_94_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_94_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_94_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_94_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_94_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_94_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_94_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_94_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_94_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_94_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_94_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_94_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_94_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_94_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_94_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_94_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_94_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_94_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_94_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_94_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_94_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_94_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_94_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_94_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_94_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_95 ( // @[mac.scala 29:63]
    .clock(PECross_95_clock),
    .reset(PECross_95_reset),
    .multiply_io_input_io_sumIn_ready(PECross_95_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_95_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_95_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_95_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_95_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_95_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_95_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_95_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_95_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_95_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_95_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_95_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_95_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_95_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_95_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_95_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_95_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_95_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_95_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_95_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_95_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_95_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_95_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_95_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_95_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_95_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_95_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_96 ( // @[mac.scala 29:63]
    .clock(PECross_96_clock),
    .reset(PECross_96_reset),
    .multiply_io_input_io_sumIn_ready(PECross_96_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_96_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_96_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_96_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_96_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_96_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_96_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_96_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_96_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_96_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_96_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_96_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_96_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_96_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_96_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_96_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_96_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_96_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_96_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_96_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_96_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_96_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_96_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_96_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_96_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_96_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_96_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_97 ( // @[mac.scala 29:63]
    .clock(PECross_97_clock),
    .reset(PECross_97_reset),
    .multiply_io_input_io_sumIn_ready(PECross_97_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_97_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_97_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_97_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_97_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_97_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_97_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_97_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_97_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_97_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_97_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_97_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_97_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_97_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_97_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_97_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_97_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_97_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_97_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_97_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_97_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_97_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_97_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_97_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_97_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_97_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_97_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_98 ( // @[mac.scala 29:63]
    .clock(PECross_98_clock),
    .reset(PECross_98_reset),
    .multiply_io_input_io_sumIn_ready(PECross_98_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_98_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_98_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_98_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_98_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_98_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_98_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_98_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_98_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_98_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_98_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_98_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_98_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_98_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_98_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_98_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_98_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_98_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_98_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_98_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_98_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_98_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_98_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_98_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_98_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_98_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_98_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_99 ( // @[mac.scala 29:63]
    .clock(PECross_99_clock),
    .reset(PECross_99_reset),
    .multiply_io_input_io_sumIn_ready(PECross_99_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_99_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_99_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_99_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_99_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_99_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_99_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_99_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_99_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_99_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_99_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_99_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_99_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_99_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_99_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_99_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_99_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_99_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_99_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_99_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_99_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_99_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_99_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_99_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_99_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_99_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_99_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_100 ( // @[mac.scala 29:63]
    .clock(PECross_100_clock),
    .reset(PECross_100_reset),
    .multiply_io_input_io_sumIn_ready(PECross_100_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_100_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_100_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_100_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_100_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_100_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_100_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_100_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_100_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_100_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_100_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_100_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_100_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_100_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_100_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_100_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_100_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_100_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_100_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_100_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_100_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_100_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_100_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_100_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_100_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_100_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_100_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_101 ( // @[mac.scala 29:63]
    .clock(PECross_101_clock),
    .reset(PECross_101_reset),
    .multiply_io_input_io_sumIn_ready(PECross_101_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_101_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_101_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_101_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_101_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_101_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_101_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_101_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_101_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_101_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_101_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_101_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_101_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_101_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_101_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_101_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_101_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_101_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_101_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_101_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_101_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_101_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_101_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_101_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_101_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_101_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_101_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_102 ( // @[mac.scala 29:63]
    .clock(PECross_102_clock),
    .reset(PECross_102_reset),
    .multiply_io_input_io_sumIn_ready(PECross_102_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_102_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_102_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_102_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_102_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_102_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_102_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_102_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_102_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_102_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_102_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_102_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_102_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_102_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_102_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_102_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_102_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_102_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_102_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_102_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_102_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_102_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_102_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_102_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_102_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_102_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_102_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_103 ( // @[mac.scala 29:63]
    .clock(PECross_103_clock),
    .reset(PECross_103_reset),
    .multiply_io_input_io_sumIn_ready(PECross_103_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_103_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_103_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_103_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_103_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_103_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_103_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_103_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_103_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_103_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_103_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_103_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_103_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_103_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_103_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_103_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_103_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_103_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_103_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_103_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_103_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_103_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_103_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_103_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_103_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_103_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_103_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_104 ( // @[mac.scala 29:63]
    .clock(PECross_104_clock),
    .reset(PECross_104_reset),
    .multiply_io_input_io_sumIn_ready(PECross_104_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_104_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_104_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_104_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_104_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_104_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_104_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_104_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_104_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_104_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_104_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_104_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_104_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_104_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_104_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_104_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_104_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_104_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_104_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_104_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_104_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_104_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_104_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_104_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_104_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_104_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_104_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_105 ( // @[mac.scala 29:63]
    .clock(PECross_105_clock),
    .reset(PECross_105_reset),
    .multiply_io_input_io_sumIn_ready(PECross_105_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_105_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_105_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_105_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_105_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_105_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_105_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_105_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_105_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_105_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_105_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_105_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_105_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_105_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_105_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_105_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_105_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_105_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_105_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_105_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_105_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_105_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_105_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_105_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_105_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_105_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_105_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_106 ( // @[mac.scala 29:63]
    .clock(PECross_106_clock),
    .reset(PECross_106_reset),
    .multiply_io_input_io_sumIn_ready(PECross_106_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_106_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_106_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_106_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_106_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_106_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_106_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_106_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_106_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_106_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_106_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_106_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_106_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_106_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_106_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_106_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_106_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_106_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_106_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_106_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_106_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_106_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_106_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_106_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_106_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_106_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_106_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_107 ( // @[mac.scala 29:63]
    .clock(PECross_107_clock),
    .reset(PECross_107_reset),
    .multiply_io_input_io_sumIn_ready(PECross_107_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_107_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_107_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_107_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_107_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_107_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_107_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_107_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_107_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_107_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_107_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_107_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_107_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_107_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_107_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_107_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_107_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_107_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_107_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_107_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_107_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_107_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_107_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_107_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_107_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_107_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_107_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_108 ( // @[mac.scala 29:63]
    .clock(PECross_108_clock),
    .reset(PECross_108_reset),
    .multiply_io_input_io_sumIn_ready(PECross_108_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_108_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_108_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_108_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_108_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_108_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_108_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_108_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_108_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_108_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_108_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_108_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_108_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_108_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_108_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_108_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_108_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_108_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_108_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_108_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_108_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_108_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_108_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_108_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_108_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_108_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_108_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_109 ( // @[mac.scala 29:63]
    .clock(PECross_109_clock),
    .reset(PECross_109_reset),
    .multiply_io_input_io_sumIn_ready(PECross_109_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_109_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_109_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_109_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_109_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_109_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_109_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_109_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_109_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_109_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_109_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_109_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_109_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_109_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_109_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_109_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_109_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_109_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_109_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_109_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_109_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_109_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_109_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_109_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_109_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_109_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_109_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_110 ( // @[mac.scala 29:63]
    .clock(PECross_110_clock),
    .reset(PECross_110_reset),
    .multiply_io_input_io_sumIn_ready(PECross_110_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_110_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_110_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_110_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_110_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_110_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_110_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_110_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_110_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_110_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_110_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_110_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_110_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_110_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_110_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_110_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_110_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_110_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_110_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_110_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_110_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_110_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_110_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_110_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_110_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_110_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_110_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_111 ( // @[mac.scala 29:63]
    .clock(PECross_111_clock),
    .reset(PECross_111_reset),
    .multiply_io_input_io_sumIn_ready(PECross_111_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_111_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_111_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_111_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_111_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_111_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_111_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_111_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_111_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_111_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_111_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_111_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_111_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_111_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_111_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_111_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_111_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_111_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_111_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_111_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_111_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_111_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_111_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_111_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_111_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_111_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_111_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_112 ( // @[mac.scala 29:63]
    .clock(PECross_112_clock),
    .reset(PECross_112_reset),
    .multiply_io_input_io_sumIn_ready(PECross_112_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_112_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_112_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_112_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_112_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_112_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_112_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_112_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_112_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_112_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_112_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_112_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_112_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_112_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_112_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_112_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_112_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_112_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_112_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_112_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_112_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_112_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_112_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_112_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_112_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_112_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_112_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_113 ( // @[mac.scala 29:63]
    .clock(PECross_113_clock),
    .reset(PECross_113_reset),
    .multiply_io_input_io_sumIn_ready(PECross_113_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_113_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_113_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_113_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_113_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_113_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_113_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_113_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_113_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_113_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_113_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_113_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_113_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_113_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_113_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_113_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_113_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_113_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_113_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_113_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_113_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_113_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_113_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_113_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_113_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_113_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_113_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_114 ( // @[mac.scala 29:63]
    .clock(PECross_114_clock),
    .reset(PECross_114_reset),
    .multiply_io_input_io_sumIn_ready(PECross_114_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_114_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_114_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_114_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_114_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_114_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_114_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_114_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_114_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_114_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_114_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_114_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_114_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_114_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_114_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_114_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_114_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_114_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_114_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_114_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_114_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_114_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_114_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_114_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_114_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_114_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_114_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_115 ( // @[mac.scala 29:63]
    .clock(PECross_115_clock),
    .reset(PECross_115_reset),
    .multiply_io_input_io_sumIn_ready(PECross_115_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_115_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_115_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_115_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_115_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_115_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_115_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_115_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_115_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_115_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_115_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_115_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_115_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_115_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_115_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_115_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_115_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_115_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_115_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_115_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_115_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_115_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_115_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_115_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_115_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_115_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_115_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_116 ( // @[mac.scala 29:63]
    .clock(PECross_116_clock),
    .reset(PECross_116_reset),
    .multiply_io_input_io_sumIn_ready(PECross_116_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_116_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_116_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_116_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_116_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_116_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_116_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_116_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_116_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_116_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_116_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_116_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_116_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_116_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_116_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_116_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_116_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_116_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_116_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_116_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_116_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_116_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_116_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_116_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_116_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_116_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_116_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_117 ( // @[mac.scala 29:63]
    .clock(PECross_117_clock),
    .reset(PECross_117_reset),
    .multiply_io_input_io_sumIn_ready(PECross_117_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_117_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_117_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_117_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_117_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_117_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_117_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_117_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_117_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_117_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_117_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_117_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_117_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_117_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_117_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_117_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_117_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_117_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_117_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_117_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_117_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_117_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_117_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_117_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_117_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_117_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_117_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_118 ( // @[mac.scala 29:63]
    .clock(PECross_118_clock),
    .reset(PECross_118_reset),
    .multiply_io_input_io_sumIn_ready(PECross_118_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_118_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_118_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_118_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_118_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_118_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_118_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_118_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_118_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_118_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_118_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_118_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_118_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_118_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_118_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_118_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_118_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_118_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_118_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_118_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_118_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_118_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_118_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_118_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_118_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_118_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_118_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_119 ( // @[mac.scala 29:63]
    .clock(PECross_119_clock),
    .reset(PECross_119_reset),
    .multiply_io_input_io_sumIn_ready(PECross_119_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_119_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_119_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_119_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_119_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_119_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_119_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_119_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_119_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_119_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_119_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_119_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_119_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_119_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_119_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_119_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_119_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_119_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_119_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_119_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_119_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_119_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_119_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_119_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_119_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_119_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_119_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_120 ( // @[mac.scala 29:63]
    .clock(PECross_120_clock),
    .reset(PECross_120_reset),
    .multiply_io_input_io_sumIn_ready(PECross_120_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_120_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_120_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_120_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_120_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_120_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_120_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_120_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_120_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_120_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_120_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_120_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_120_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_120_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_120_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_120_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_120_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_120_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_120_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_120_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_120_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_120_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_120_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_120_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_120_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_120_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_120_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_121 ( // @[mac.scala 29:63]
    .clock(PECross_121_clock),
    .reset(PECross_121_reset),
    .multiply_io_input_io_sumIn_ready(PECross_121_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_121_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_121_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_121_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_121_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_121_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_121_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_121_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_121_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_121_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_121_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_121_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_121_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_121_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_121_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_121_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_121_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_121_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_121_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_121_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_121_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_121_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_121_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_121_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_121_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_121_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_121_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_122 ( // @[mac.scala 29:63]
    .clock(PECross_122_clock),
    .reset(PECross_122_reset),
    .multiply_io_input_io_sumIn_ready(PECross_122_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_122_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_122_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_122_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_122_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_122_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_122_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_122_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_122_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_122_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_122_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_122_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_122_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_122_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_122_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_122_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_122_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_122_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_122_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_122_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_122_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_122_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_122_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_122_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_122_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_122_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_122_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_123 ( // @[mac.scala 29:63]
    .clock(PECross_123_clock),
    .reset(PECross_123_reset),
    .multiply_io_input_io_sumIn_ready(PECross_123_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_123_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_123_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_123_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_123_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_123_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_123_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_123_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_123_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_123_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_123_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_123_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_123_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_123_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_123_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_123_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_123_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_123_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_123_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_123_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_123_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_123_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_123_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_123_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_123_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_123_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_123_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_124 ( // @[mac.scala 29:63]
    .clock(PECross_124_clock),
    .reset(PECross_124_reset),
    .multiply_io_input_io_sumIn_ready(PECross_124_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_124_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_124_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_124_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_124_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_124_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_124_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_124_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_124_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_124_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_124_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_124_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_124_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_124_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_124_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_124_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_124_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_124_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_124_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_124_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_124_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_124_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_124_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_124_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_124_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_124_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_124_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_125 ( // @[mac.scala 29:63]
    .clock(PECross_125_clock),
    .reset(PECross_125_reset),
    .multiply_io_input_io_sumIn_ready(PECross_125_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_125_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_125_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_125_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_125_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_125_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_125_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_125_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_125_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_125_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_125_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_125_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_125_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_125_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_125_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_125_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_125_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_125_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_125_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_125_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_125_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_125_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_125_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_125_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_125_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_125_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_125_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_126 ( // @[mac.scala 29:63]
    .clock(PECross_126_clock),
    .reset(PECross_126_reset),
    .multiply_io_input_io_sumIn_ready(PECross_126_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_126_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_126_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_126_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_126_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_126_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_126_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_126_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_126_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_126_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_126_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_126_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_126_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_126_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_126_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_126_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_126_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_126_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_126_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_126_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_126_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_126_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_126_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_126_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_126_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_126_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_126_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_127 ( // @[mac.scala 29:63]
    .clock(PECross_127_clock),
    .reset(PECross_127_reset),
    .multiply_io_input_io_sumIn_ready(PECross_127_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_127_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_127_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_127_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_127_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_127_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_127_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_127_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_127_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_127_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_127_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_127_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_127_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_127_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_127_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_127_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_127_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_127_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_127_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_127_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_127_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_127_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_127_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_127_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_127_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_127_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_127_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_128 ( // @[mac.scala 29:63]
    .clock(PECross_128_clock),
    .reset(PECross_128_reset),
    .multiply_io_input_io_sumIn_ready(PECross_128_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_128_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_128_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_128_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_128_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_128_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_128_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_128_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_128_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_128_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_128_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_128_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_128_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_128_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_128_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_128_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_128_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_128_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_128_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_128_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_128_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_128_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_128_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_128_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_128_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_128_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_128_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_129 ( // @[mac.scala 29:63]
    .clock(PECross_129_clock),
    .reset(PECross_129_reset),
    .multiply_io_input_io_sumIn_ready(PECross_129_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_129_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_129_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_129_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_129_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_129_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_129_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_129_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_129_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_129_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_129_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_129_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_129_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_129_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_129_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_129_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_129_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_129_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_129_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_129_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_129_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_129_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_129_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_129_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_129_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_129_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_129_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_130 ( // @[mac.scala 29:63]
    .clock(PECross_130_clock),
    .reset(PECross_130_reset),
    .multiply_io_input_io_sumIn_ready(PECross_130_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_130_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_130_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_130_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_130_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_130_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_130_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_130_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_130_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_130_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_130_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_130_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_130_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_130_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_130_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_130_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_130_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_130_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_130_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_130_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_130_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_130_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_130_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_130_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_130_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_130_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_130_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_131 ( // @[mac.scala 29:63]
    .clock(PECross_131_clock),
    .reset(PECross_131_reset),
    .multiply_io_input_io_sumIn_ready(PECross_131_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_131_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_131_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_131_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_131_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_131_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_131_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_131_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_131_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_131_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_131_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_131_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_131_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_131_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_131_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_131_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_131_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_131_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_131_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_131_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_131_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_131_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_131_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_131_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_131_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_131_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_131_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_132 ( // @[mac.scala 29:63]
    .clock(PECross_132_clock),
    .reset(PECross_132_reset),
    .multiply_io_input_io_sumIn_ready(PECross_132_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_132_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_132_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_132_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_132_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_132_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_132_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_132_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_132_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_132_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_132_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_132_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_132_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_132_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_132_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_132_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_132_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_132_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_132_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_132_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_132_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_132_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_132_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_132_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_132_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_132_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_132_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_133 ( // @[mac.scala 29:63]
    .clock(PECross_133_clock),
    .reset(PECross_133_reset),
    .multiply_io_input_io_sumIn_ready(PECross_133_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_133_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_133_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_133_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_133_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_133_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_133_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_133_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_133_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_133_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_133_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_133_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_133_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_133_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_133_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_133_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_133_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_133_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_133_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_133_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_133_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_133_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_133_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_133_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_133_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_133_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_133_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_134 ( // @[mac.scala 29:63]
    .clock(PECross_134_clock),
    .reset(PECross_134_reset),
    .multiply_io_input_io_sumIn_ready(PECross_134_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_134_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_134_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_134_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_134_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_134_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_134_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_134_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_134_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_134_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_134_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_134_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_134_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_134_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_134_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_134_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_134_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_134_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_134_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_134_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_134_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_134_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_134_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_134_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_134_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_134_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_134_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_135 ( // @[mac.scala 29:63]
    .clock(PECross_135_clock),
    .reset(PECross_135_reset),
    .multiply_io_input_io_sumIn_ready(PECross_135_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_135_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_135_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_135_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_135_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_135_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_135_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_135_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_135_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_135_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_135_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_135_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_135_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_135_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_135_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_135_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_135_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_135_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_135_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_135_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_135_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_135_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_135_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_135_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_135_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_135_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_135_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_136 ( // @[mac.scala 29:63]
    .clock(PECross_136_clock),
    .reset(PECross_136_reset),
    .multiply_io_input_io_sumIn_ready(PECross_136_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_136_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_136_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_136_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_136_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_136_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_136_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_136_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_136_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_136_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_136_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_136_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_136_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_136_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_136_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_136_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_136_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_136_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_136_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_136_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_136_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_136_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_136_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_136_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_136_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_136_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_136_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_137 ( // @[mac.scala 29:63]
    .clock(PECross_137_clock),
    .reset(PECross_137_reset),
    .multiply_io_input_io_sumIn_ready(PECross_137_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_137_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_137_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_137_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_137_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_137_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_137_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_137_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_137_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_137_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_137_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_137_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_137_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_137_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_137_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_137_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_137_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_137_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_137_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_137_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_137_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_137_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_137_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_137_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_137_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_137_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_137_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_138 ( // @[mac.scala 29:63]
    .clock(PECross_138_clock),
    .reset(PECross_138_reset),
    .multiply_io_input_io_sumIn_ready(PECross_138_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_138_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_138_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_138_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_138_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_138_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_138_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_138_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_138_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_138_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_138_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_138_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_138_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_138_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_138_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_138_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_138_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_138_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_138_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_138_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_138_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_138_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_138_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_138_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_138_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_138_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_138_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_139 ( // @[mac.scala 29:63]
    .clock(PECross_139_clock),
    .reset(PECross_139_reset),
    .multiply_io_input_io_sumIn_ready(PECross_139_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_139_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_139_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_139_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_139_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_139_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_139_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_139_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_139_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_139_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_139_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_139_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_139_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_139_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_139_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_139_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_139_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_139_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_139_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_139_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_139_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_139_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_139_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_139_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_139_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_139_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_139_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_140 ( // @[mac.scala 29:63]
    .clock(PECross_140_clock),
    .reset(PECross_140_reset),
    .multiply_io_input_io_sumIn_ready(PECross_140_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_140_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_140_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_140_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_140_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_140_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_140_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_140_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_140_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_140_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_140_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_140_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_140_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_140_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_140_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_140_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_140_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_140_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_140_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_140_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_140_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_140_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_140_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_140_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_140_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_140_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_140_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_141 ( // @[mac.scala 29:63]
    .clock(PECross_141_clock),
    .reset(PECross_141_reset),
    .multiply_io_input_io_sumIn_ready(PECross_141_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_141_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_141_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_141_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_141_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_141_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_141_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_141_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_141_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_141_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_141_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_141_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_141_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_141_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_141_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_141_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_141_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_141_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_141_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_141_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_141_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_141_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_141_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_141_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_141_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_141_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_141_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_142 ( // @[mac.scala 29:63]
    .clock(PECross_142_clock),
    .reset(PECross_142_reset),
    .multiply_io_input_io_sumIn_ready(PECross_142_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_142_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_142_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_142_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_142_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_142_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_142_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_142_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_142_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_142_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_142_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_142_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_142_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_142_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_142_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_142_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_142_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_142_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_142_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_142_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_142_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_142_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_142_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_142_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_142_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_142_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_142_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_143 ( // @[mac.scala 29:63]
    .clock(PECross_143_clock),
    .reset(PECross_143_reset),
    .multiply_io_input_io_sumIn_ready(PECross_143_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_143_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_143_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_143_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_143_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_143_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_143_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_143_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_143_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_143_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_143_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_143_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_143_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_143_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_143_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_143_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_143_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_143_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_143_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_143_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_143_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_143_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_143_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_143_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_143_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_143_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_143_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_144 ( // @[mac.scala 29:63]
    .clock(PECross_144_clock),
    .reset(PECross_144_reset),
    .multiply_io_input_io_sumIn_ready(PECross_144_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_144_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_144_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_144_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_144_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_144_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_144_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_144_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_144_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_144_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_144_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_144_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_144_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_144_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_144_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_144_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_144_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_144_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_144_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_144_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_144_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_144_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_144_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_144_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_144_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_144_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_144_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_145 ( // @[mac.scala 29:63]
    .clock(PECross_145_clock),
    .reset(PECross_145_reset),
    .multiply_io_input_io_sumIn_ready(PECross_145_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_145_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_145_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_145_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_145_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_145_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_145_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_145_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_145_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_145_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_145_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_145_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_145_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_145_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_145_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_145_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_145_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_145_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_145_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_145_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_145_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_145_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_145_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_145_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_145_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_145_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_145_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_146 ( // @[mac.scala 29:63]
    .clock(PECross_146_clock),
    .reset(PECross_146_reset),
    .multiply_io_input_io_sumIn_ready(PECross_146_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_146_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_146_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_146_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_146_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_146_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_146_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_146_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_146_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_146_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_146_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_146_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_146_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_146_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_146_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_146_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_146_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_146_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_146_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_146_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_146_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_146_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_146_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_146_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_146_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_146_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_146_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_147 ( // @[mac.scala 29:63]
    .clock(PECross_147_clock),
    .reset(PECross_147_reset),
    .multiply_io_input_io_sumIn_ready(PECross_147_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_147_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_147_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_147_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_147_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_147_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_147_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_147_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_147_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_147_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_147_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_147_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_147_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_147_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_147_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_147_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_147_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_147_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_147_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_147_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_147_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_147_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_147_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_147_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_147_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_147_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_147_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_148 ( // @[mac.scala 29:63]
    .clock(PECross_148_clock),
    .reset(PECross_148_reset),
    .multiply_io_input_io_sumIn_ready(PECross_148_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_148_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_148_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_148_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_148_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_148_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_148_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_148_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_148_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_148_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_148_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_148_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_148_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_148_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_148_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_148_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_148_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_148_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_148_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_148_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_148_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_148_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_148_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_148_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_148_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_148_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_148_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_149 ( // @[mac.scala 29:63]
    .clock(PECross_149_clock),
    .reset(PECross_149_reset),
    .multiply_io_input_io_sumIn_ready(PECross_149_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_149_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_149_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_149_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_149_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_149_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_149_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_149_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_149_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_149_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_149_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_149_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_149_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_149_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_149_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_149_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_149_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_149_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_149_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_149_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_149_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_149_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_149_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_149_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_149_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_149_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_149_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_150 ( // @[mac.scala 29:63]
    .clock(PECross_150_clock),
    .reset(PECross_150_reset),
    .multiply_io_input_io_sumIn_ready(PECross_150_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_150_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_150_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_150_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_150_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_150_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_150_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_150_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_150_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_150_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_150_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_150_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_150_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_150_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_150_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_150_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_150_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_150_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_150_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_150_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_150_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_150_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_150_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_150_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_150_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_150_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_150_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_151 ( // @[mac.scala 29:63]
    .clock(PECross_151_clock),
    .reset(PECross_151_reset),
    .multiply_io_input_io_sumIn_ready(PECross_151_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_151_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_151_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_151_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_151_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_151_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_151_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_151_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_151_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_151_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_151_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_151_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_151_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_151_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_151_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_151_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_151_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_151_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_151_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_151_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_151_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_151_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_151_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_151_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_151_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_151_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_151_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_152 ( // @[mac.scala 29:63]
    .clock(PECross_152_clock),
    .reset(PECross_152_reset),
    .multiply_io_input_io_sumIn_ready(PECross_152_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_152_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_152_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_152_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_152_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_152_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_152_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_152_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_152_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_152_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_152_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_152_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_152_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_152_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_152_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_152_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_152_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_152_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_152_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_152_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_152_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_152_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_152_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_152_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_152_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_152_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_152_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_153 ( // @[mac.scala 29:63]
    .clock(PECross_153_clock),
    .reset(PECross_153_reset),
    .multiply_io_input_io_sumIn_ready(PECross_153_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_153_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_153_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_153_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_153_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_153_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_153_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_153_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_153_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_153_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_153_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_153_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_153_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_153_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_153_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_153_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_153_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_153_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_153_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_153_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_153_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_153_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_153_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_153_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_153_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_153_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_153_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_154 ( // @[mac.scala 29:63]
    .clock(PECross_154_clock),
    .reset(PECross_154_reset),
    .multiply_io_input_io_sumIn_ready(PECross_154_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_154_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_154_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_154_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_154_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_154_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_154_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_154_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_154_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_154_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_154_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_154_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_154_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_154_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_154_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_154_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_154_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_154_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_154_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_154_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_154_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_154_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_154_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_154_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_154_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_154_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_154_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_155 ( // @[mac.scala 29:63]
    .clock(PECross_155_clock),
    .reset(PECross_155_reset),
    .multiply_io_input_io_sumIn_ready(PECross_155_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_155_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_155_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_155_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_155_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_155_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_155_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_155_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_155_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_155_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_155_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_155_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_155_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_155_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_155_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_155_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_155_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_155_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_155_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_155_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_155_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_155_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_155_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_155_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_155_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_155_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_155_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_156 ( // @[mac.scala 29:63]
    .clock(PECross_156_clock),
    .reset(PECross_156_reset),
    .multiply_io_input_io_sumIn_ready(PECross_156_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_156_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_156_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_156_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_156_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_156_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_156_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_156_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_156_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_156_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_156_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_156_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_156_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_156_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_156_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_156_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_156_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_156_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_156_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_156_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_156_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_156_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_156_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_156_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_156_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_156_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_156_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_157 ( // @[mac.scala 29:63]
    .clock(PECross_157_clock),
    .reset(PECross_157_reset),
    .multiply_io_input_io_sumIn_ready(PECross_157_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_157_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_157_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_157_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_157_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_157_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_157_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_157_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_157_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_157_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_157_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_157_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_157_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_157_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_157_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_157_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_157_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_157_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_157_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_157_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_157_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_157_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_157_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_157_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_157_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_157_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_157_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_158 ( // @[mac.scala 29:63]
    .clock(PECross_158_clock),
    .reset(PECross_158_reset),
    .multiply_io_input_io_sumIn_ready(PECross_158_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_158_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_158_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_158_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_158_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_158_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_158_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_158_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_158_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_158_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_158_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_158_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_158_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_158_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_158_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_158_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_158_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_158_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_158_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_158_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_158_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_158_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_158_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_158_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_158_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_158_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_158_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_159 ( // @[mac.scala 29:63]
    .clock(PECross_159_clock),
    .reset(PECross_159_reset),
    .multiply_io_input_io_sumIn_ready(PECross_159_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_159_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_159_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_159_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_159_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_159_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_159_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_159_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_159_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_159_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_159_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_159_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_159_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_159_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_159_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_159_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_159_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_159_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_159_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_159_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_159_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_159_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_159_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_159_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_159_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_159_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_159_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_160 ( // @[mac.scala 29:63]
    .clock(PECross_160_clock),
    .reset(PECross_160_reset),
    .multiply_io_input_io_sumIn_ready(PECross_160_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_160_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_160_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_160_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_160_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_160_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_160_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_160_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_160_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_160_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_160_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_160_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_160_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_160_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_160_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_160_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_160_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_160_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_160_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_160_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_160_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_160_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_160_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_160_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_160_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_160_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_160_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_161 ( // @[mac.scala 29:63]
    .clock(PECross_161_clock),
    .reset(PECross_161_reset),
    .multiply_io_input_io_sumIn_ready(PECross_161_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_161_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_161_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_161_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_161_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_161_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_161_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_161_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_161_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_161_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_161_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_161_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_161_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_161_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_161_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_161_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_161_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_161_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_161_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_161_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_161_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_161_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_161_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_161_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_161_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_161_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_161_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_162 ( // @[mac.scala 29:63]
    .clock(PECross_162_clock),
    .reset(PECross_162_reset),
    .multiply_io_input_io_sumIn_ready(PECross_162_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_162_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_162_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_162_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_162_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_162_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_162_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_162_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_162_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_162_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_162_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_162_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_162_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_162_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_162_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_162_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_162_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_162_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_162_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_162_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_162_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_162_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_162_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_162_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_162_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_162_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_162_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_163 ( // @[mac.scala 29:63]
    .clock(PECross_163_clock),
    .reset(PECross_163_reset),
    .multiply_io_input_io_sumIn_ready(PECross_163_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_163_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_163_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_163_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_163_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_163_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_163_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_163_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_163_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_163_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_163_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_163_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_163_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_163_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_163_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_163_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_163_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_163_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_163_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_163_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_163_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_163_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_163_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_163_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_163_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_163_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_163_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_164 ( // @[mac.scala 29:63]
    .clock(PECross_164_clock),
    .reset(PECross_164_reset),
    .multiply_io_input_io_sumIn_ready(PECross_164_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_164_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_164_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_164_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_164_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_164_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_164_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_164_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_164_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_164_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_164_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_164_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_164_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_164_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_164_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_164_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_164_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_164_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_164_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_164_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_164_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_164_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_164_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_164_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_164_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_164_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_164_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_165 ( // @[mac.scala 29:63]
    .clock(PECross_165_clock),
    .reset(PECross_165_reset),
    .multiply_io_input_io_sumIn_ready(PECross_165_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_165_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_165_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_165_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_165_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_165_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_165_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_165_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_165_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_165_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_165_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_165_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_165_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_165_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_165_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_165_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_165_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_165_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_165_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_165_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_165_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_165_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_165_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_165_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_165_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_165_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_165_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_166 ( // @[mac.scala 29:63]
    .clock(PECross_166_clock),
    .reset(PECross_166_reset),
    .multiply_io_input_io_sumIn_ready(PECross_166_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_166_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_166_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_166_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_166_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_166_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_166_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_166_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_166_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_166_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_166_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_166_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_166_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_166_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_166_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_166_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_166_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_166_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_166_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_166_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_166_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_166_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_166_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_166_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_166_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_166_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_166_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_167 ( // @[mac.scala 29:63]
    .clock(PECross_167_clock),
    .reset(PECross_167_reset),
    .multiply_io_input_io_sumIn_ready(PECross_167_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_167_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_167_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_167_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_167_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_167_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_167_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_167_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_167_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_167_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_167_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_167_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_167_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_167_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_167_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_167_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_167_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_167_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_167_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_167_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_167_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_167_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_167_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_167_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_167_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_167_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_167_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_168 ( // @[mac.scala 29:63]
    .clock(PECross_168_clock),
    .reset(PECross_168_reset),
    .multiply_io_input_io_sumIn_ready(PECross_168_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_168_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_168_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_168_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_168_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_168_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_168_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_168_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_168_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_168_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_168_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_168_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_168_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_168_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_168_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_168_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_168_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_168_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_168_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_168_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_168_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_168_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_168_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_168_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_168_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_168_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_168_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_169 ( // @[mac.scala 29:63]
    .clock(PECross_169_clock),
    .reset(PECross_169_reset),
    .multiply_io_input_io_sumIn_ready(PECross_169_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_169_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_169_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_169_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_169_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_169_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_169_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_169_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_169_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_169_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_169_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_169_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_169_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_169_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_169_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_169_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_169_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_169_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_169_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_169_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_169_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_169_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_169_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_169_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_169_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_169_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_169_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_170 ( // @[mac.scala 29:63]
    .clock(PECross_170_clock),
    .reset(PECross_170_reset),
    .multiply_io_input_io_sumIn_ready(PECross_170_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_170_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_170_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_170_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_170_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_170_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_170_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_170_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_170_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_170_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_170_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_170_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_170_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_170_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_170_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_170_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_170_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_170_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_170_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_170_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_170_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_170_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_170_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_170_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_170_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_170_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_170_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_171 ( // @[mac.scala 29:63]
    .clock(PECross_171_clock),
    .reset(PECross_171_reset),
    .multiply_io_input_io_sumIn_ready(PECross_171_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_171_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_171_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_171_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_171_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_171_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_171_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_171_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_171_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_171_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_171_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_171_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_171_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_171_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_171_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_171_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_171_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_171_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_171_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_171_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_171_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_171_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_171_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_171_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_171_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_171_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_171_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_172 ( // @[mac.scala 29:63]
    .clock(PECross_172_clock),
    .reset(PECross_172_reset),
    .multiply_io_input_io_sumIn_ready(PECross_172_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_172_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_172_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_172_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_172_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_172_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_172_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_172_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_172_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_172_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_172_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_172_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_172_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_172_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_172_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_172_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_172_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_172_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_172_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_172_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_172_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_172_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_172_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_172_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_172_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_172_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_172_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_173 ( // @[mac.scala 29:63]
    .clock(PECross_173_clock),
    .reset(PECross_173_reset),
    .multiply_io_input_io_sumIn_ready(PECross_173_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_173_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_173_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_173_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_173_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_173_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_173_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_173_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_173_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_173_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_173_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_173_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_173_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_173_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_173_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_173_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_173_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_173_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_173_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_173_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_173_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_173_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_173_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_173_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_173_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_173_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_173_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_174 ( // @[mac.scala 29:63]
    .clock(PECross_174_clock),
    .reset(PECross_174_reset),
    .multiply_io_input_io_sumIn_ready(PECross_174_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_174_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_174_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_174_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_174_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_174_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_174_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_174_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_174_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_174_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_174_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_174_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_174_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_174_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_174_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_174_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_174_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_174_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_174_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_174_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_174_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_174_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_174_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_174_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_174_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_174_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_174_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_175 ( // @[mac.scala 29:63]
    .clock(PECross_175_clock),
    .reset(PECross_175_reset),
    .multiply_io_input_io_sumIn_ready(PECross_175_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_175_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_175_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_175_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_175_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_175_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_175_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_175_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_175_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_175_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_175_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_175_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_175_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_175_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_175_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_175_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_175_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_175_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_175_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_175_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_175_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_175_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_175_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_175_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_175_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_175_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_175_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_176 ( // @[mac.scala 29:63]
    .clock(PECross_176_clock),
    .reset(PECross_176_reset),
    .multiply_io_input_io_sumIn_ready(PECross_176_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_176_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_176_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_176_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_176_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_176_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_176_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_176_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_176_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_176_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_176_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_176_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_176_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_176_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_176_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_176_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_176_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_176_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_176_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_176_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_176_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_176_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_176_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_176_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_176_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_176_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_176_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_177 ( // @[mac.scala 29:63]
    .clock(PECross_177_clock),
    .reset(PECross_177_reset),
    .multiply_io_input_io_sumIn_ready(PECross_177_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_177_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_177_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_177_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_177_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_177_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_177_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_177_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_177_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_177_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_177_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_177_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_177_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_177_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_177_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_177_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_177_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_177_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_177_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_177_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_177_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_177_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_177_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_177_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_177_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_177_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_177_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_178 ( // @[mac.scala 29:63]
    .clock(PECross_178_clock),
    .reset(PECross_178_reset),
    .multiply_io_input_io_sumIn_ready(PECross_178_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_178_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_178_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_178_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_178_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_178_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_178_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_178_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_178_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_178_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_178_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_178_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_178_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_178_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_178_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_178_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_178_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_178_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_178_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_178_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_178_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_178_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_178_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_178_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_178_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_178_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_178_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_179 ( // @[mac.scala 29:63]
    .clock(PECross_179_clock),
    .reset(PECross_179_reset),
    .multiply_io_input_io_sumIn_ready(PECross_179_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_179_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_179_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_179_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_179_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_179_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_179_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_179_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_179_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_179_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_179_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_179_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_179_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_179_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_179_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_179_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_179_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_179_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_179_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_179_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_179_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_179_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_179_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_179_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_179_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_179_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_179_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_180 ( // @[mac.scala 29:63]
    .clock(PECross_180_clock),
    .reset(PECross_180_reset),
    .multiply_io_input_io_sumIn_ready(PECross_180_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_180_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_180_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_180_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_180_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_180_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_180_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_180_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_180_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_180_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_180_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_180_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_180_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_180_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_180_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_180_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_180_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_180_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_180_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_180_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_180_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_180_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_180_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_180_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_180_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_180_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_180_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_181 ( // @[mac.scala 29:63]
    .clock(PECross_181_clock),
    .reset(PECross_181_reset),
    .multiply_io_input_io_sumIn_ready(PECross_181_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_181_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_181_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_181_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_181_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_181_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_181_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_181_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_181_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_181_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_181_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_181_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_181_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_181_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_181_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_181_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_181_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_181_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_181_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_181_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_181_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_181_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_181_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_181_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_181_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_181_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_181_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_182 ( // @[mac.scala 29:63]
    .clock(PECross_182_clock),
    .reset(PECross_182_reset),
    .multiply_io_input_io_sumIn_ready(PECross_182_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_182_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_182_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_182_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_182_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_182_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_182_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_182_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_182_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_182_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_182_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_182_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_182_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_182_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_182_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_182_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_182_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_182_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_182_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_182_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_182_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_182_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_182_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_182_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_182_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_182_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_182_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_183 ( // @[mac.scala 29:63]
    .clock(PECross_183_clock),
    .reset(PECross_183_reset),
    .multiply_io_input_io_sumIn_ready(PECross_183_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_183_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_183_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_183_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_183_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_183_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_183_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_183_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_183_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_183_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_183_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_183_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_183_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_183_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_183_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_183_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_183_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_183_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_183_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_183_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_183_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_183_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_183_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_183_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_183_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_183_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_183_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_184 ( // @[mac.scala 29:63]
    .clock(PECross_184_clock),
    .reset(PECross_184_reset),
    .multiply_io_input_io_sumIn_ready(PECross_184_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_184_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_184_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_184_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_184_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_184_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_184_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_184_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_184_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_184_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_184_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_184_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_184_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_184_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_184_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_184_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_184_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_184_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_184_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_184_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_184_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_184_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_184_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_184_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_184_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_184_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_184_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_185 ( // @[mac.scala 29:63]
    .clock(PECross_185_clock),
    .reset(PECross_185_reset),
    .multiply_io_input_io_sumIn_ready(PECross_185_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_185_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_185_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_185_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_185_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_185_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_185_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_185_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_185_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_185_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_185_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_185_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_185_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_185_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_185_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_185_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_185_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_185_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_185_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_185_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_185_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_185_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_185_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_185_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_185_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_185_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_185_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_186 ( // @[mac.scala 29:63]
    .clock(PECross_186_clock),
    .reset(PECross_186_reset),
    .multiply_io_input_io_sumIn_ready(PECross_186_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_186_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_186_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_186_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_186_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_186_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_186_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_186_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_186_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_186_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_186_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_186_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_186_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_186_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_186_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_186_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_186_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_186_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_186_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_186_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_186_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_186_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_186_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_186_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_186_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_186_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_186_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_187 ( // @[mac.scala 29:63]
    .clock(PECross_187_clock),
    .reset(PECross_187_reset),
    .multiply_io_input_io_sumIn_ready(PECross_187_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_187_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_187_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_187_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_187_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_187_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_187_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_187_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_187_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_187_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_187_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_187_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_187_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_187_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_187_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_187_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_187_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_187_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_187_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_187_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_187_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_187_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_187_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_187_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_187_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_187_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_187_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_188 ( // @[mac.scala 29:63]
    .clock(PECross_188_clock),
    .reset(PECross_188_reset),
    .multiply_io_input_io_sumIn_ready(PECross_188_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_188_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_188_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_188_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_188_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_188_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_188_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_188_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_188_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_188_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_188_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_188_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_188_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_188_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_188_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_188_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_188_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_188_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_188_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_188_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_188_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_188_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_188_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_188_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_188_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_188_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_188_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_189 ( // @[mac.scala 29:63]
    .clock(PECross_189_clock),
    .reset(PECross_189_reset),
    .multiply_io_input_io_sumIn_ready(PECross_189_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_189_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_189_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_189_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_189_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_189_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_189_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_189_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_189_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_189_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_189_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_189_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_189_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_189_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_189_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_189_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_189_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_189_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_189_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_189_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_189_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_189_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_189_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_189_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_189_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_189_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_189_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_190 ( // @[mac.scala 29:63]
    .clock(PECross_190_clock),
    .reset(PECross_190_reset),
    .multiply_io_input_io_sumIn_ready(PECross_190_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_190_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_190_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_190_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_190_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_190_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_190_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_190_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_190_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_190_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_190_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_190_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_190_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_190_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_190_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_190_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_190_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_190_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_190_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_190_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_190_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_190_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_190_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_190_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_190_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_190_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_190_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_191 ( // @[mac.scala 29:63]
    .clock(PECross_191_clock),
    .reset(PECross_191_reset),
    .multiply_io_input_io_sumIn_ready(PECross_191_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_191_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_191_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_191_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_191_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_191_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_191_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_191_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_191_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_191_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_191_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_191_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_191_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_191_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_191_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_191_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_191_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_191_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_191_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_191_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_191_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_191_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_191_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_191_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_191_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_191_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_191_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_192 ( // @[mac.scala 29:63]
    .clock(PECross_192_clock),
    .reset(PECross_192_reset),
    .multiply_io_input_io_sumIn_ready(PECross_192_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_192_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_192_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_192_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_192_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_192_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_192_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_192_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_192_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_192_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_192_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_192_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_192_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_192_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_192_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_192_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_192_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_192_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_192_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_192_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_192_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_192_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_192_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_192_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_192_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_192_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_192_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_193 ( // @[mac.scala 29:63]
    .clock(PECross_193_clock),
    .reset(PECross_193_reset),
    .multiply_io_input_io_sumIn_ready(PECross_193_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_193_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_193_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_193_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_193_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_193_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_193_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_193_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_193_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_193_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_193_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_193_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_193_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_193_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_193_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_193_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_193_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_193_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_193_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_193_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_193_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_193_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_193_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_193_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_193_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_193_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_193_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_194 ( // @[mac.scala 29:63]
    .clock(PECross_194_clock),
    .reset(PECross_194_reset),
    .multiply_io_input_io_sumIn_ready(PECross_194_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_194_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_194_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_194_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_194_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_194_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_194_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_194_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_194_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_194_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_194_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_194_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_194_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_194_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_194_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_194_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_194_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_194_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_194_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_194_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_194_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_194_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_194_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_194_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_194_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_194_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_194_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_195 ( // @[mac.scala 29:63]
    .clock(PECross_195_clock),
    .reset(PECross_195_reset),
    .multiply_io_input_io_sumIn_ready(PECross_195_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_195_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_195_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_195_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_195_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_195_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_195_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_195_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_195_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_195_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_195_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_195_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_195_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_195_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_195_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_195_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_195_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_195_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_195_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_195_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_195_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_195_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_195_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_195_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_195_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_195_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_195_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_196 ( // @[mac.scala 29:63]
    .clock(PECross_196_clock),
    .reset(PECross_196_reset),
    .multiply_io_input_io_sumIn_ready(PECross_196_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_196_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_196_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_196_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_196_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_196_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_196_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_196_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_196_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_196_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_196_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_196_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_196_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_196_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_196_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_196_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_196_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_196_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_196_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_196_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_196_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_196_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_196_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_196_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_196_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_196_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_196_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_197 ( // @[mac.scala 29:63]
    .clock(PECross_197_clock),
    .reset(PECross_197_reset),
    .multiply_io_input_io_sumIn_ready(PECross_197_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_197_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_197_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_197_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_197_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_197_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_197_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_197_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_197_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_197_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_197_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_197_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_197_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_197_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_197_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_197_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_197_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_197_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_197_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_197_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_197_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_197_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_197_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_197_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_197_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_197_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_197_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_198 ( // @[mac.scala 29:63]
    .clock(PECross_198_clock),
    .reset(PECross_198_reset),
    .multiply_io_input_io_sumIn_ready(PECross_198_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_198_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_198_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_198_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_198_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_198_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_198_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_198_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_198_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_198_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_198_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_198_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_198_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_198_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_198_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_198_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_198_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_198_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_198_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_198_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_198_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_198_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_198_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_198_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_198_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_198_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_198_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_199 ( // @[mac.scala 29:63]
    .clock(PECross_199_clock),
    .reset(PECross_199_reset),
    .multiply_io_input_io_sumIn_ready(PECross_199_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_199_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_199_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_199_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_199_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_199_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_199_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_199_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_199_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_199_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_199_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_199_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_199_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_199_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_199_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_199_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_199_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_199_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_199_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_199_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_199_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_199_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_199_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_199_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_199_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_199_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_199_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_200 ( // @[mac.scala 29:63]
    .clock(PECross_200_clock),
    .reset(PECross_200_reset),
    .multiply_io_input_io_sumIn_ready(PECross_200_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_200_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_200_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_200_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_200_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_200_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_200_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_200_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_200_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_200_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_200_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_200_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_200_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_200_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_200_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_200_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_200_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_200_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_200_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_200_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_200_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_200_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_200_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_200_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_200_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_200_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_200_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_201 ( // @[mac.scala 29:63]
    .clock(PECross_201_clock),
    .reset(PECross_201_reset),
    .multiply_io_input_io_sumIn_ready(PECross_201_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_201_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_201_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_201_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_201_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_201_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_201_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_201_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_201_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_201_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_201_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_201_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_201_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_201_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_201_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_201_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_201_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_201_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_201_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_201_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_201_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_201_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_201_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_201_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_201_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_201_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_201_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_202 ( // @[mac.scala 29:63]
    .clock(PECross_202_clock),
    .reset(PECross_202_reset),
    .multiply_io_input_io_sumIn_ready(PECross_202_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_202_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_202_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_202_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_202_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_202_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_202_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_202_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_202_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_202_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_202_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_202_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_202_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_202_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_202_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_202_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_202_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_202_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_202_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_202_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_202_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_202_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_202_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_202_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_202_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_202_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_202_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_203 ( // @[mac.scala 29:63]
    .clock(PECross_203_clock),
    .reset(PECross_203_reset),
    .multiply_io_input_io_sumIn_ready(PECross_203_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_203_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_203_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_203_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_203_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_203_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_203_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_203_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_203_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_203_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_203_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_203_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_203_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_203_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_203_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_203_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_203_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_203_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_203_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_203_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_203_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_203_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_203_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_203_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_203_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_203_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_203_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_204 ( // @[mac.scala 29:63]
    .clock(PECross_204_clock),
    .reset(PECross_204_reset),
    .multiply_io_input_io_sumIn_ready(PECross_204_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_204_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_204_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_204_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_204_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_204_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_204_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_204_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_204_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_204_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_204_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_204_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_204_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_204_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_204_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_204_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_204_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_204_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_204_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_204_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_204_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_204_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_204_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_204_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_204_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_204_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_204_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_205 ( // @[mac.scala 29:63]
    .clock(PECross_205_clock),
    .reset(PECross_205_reset),
    .multiply_io_input_io_sumIn_ready(PECross_205_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_205_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_205_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_205_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_205_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_205_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_205_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_205_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_205_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_205_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_205_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_205_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_205_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_205_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_205_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_205_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_205_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_205_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_205_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_205_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_205_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_205_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_205_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_205_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_205_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_205_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_205_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_206 ( // @[mac.scala 29:63]
    .clock(PECross_206_clock),
    .reset(PECross_206_reset),
    .multiply_io_input_io_sumIn_ready(PECross_206_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_206_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_206_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_206_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_206_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_206_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_206_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_206_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_206_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_206_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_206_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_206_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_206_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_206_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_206_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_206_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_206_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_206_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_206_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_206_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_206_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_206_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_206_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_206_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_206_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_206_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_206_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_207 ( // @[mac.scala 29:63]
    .clock(PECross_207_clock),
    .reset(PECross_207_reset),
    .multiply_io_input_io_sumIn_ready(PECross_207_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_207_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_207_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_207_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_207_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_207_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_207_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_207_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_207_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_207_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_207_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_207_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_207_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_207_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_207_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_207_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_207_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_207_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_207_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_207_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_207_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_207_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_207_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_207_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_207_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_207_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_207_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_208 ( // @[mac.scala 29:63]
    .clock(PECross_208_clock),
    .reset(PECross_208_reset),
    .multiply_io_input_io_sumIn_ready(PECross_208_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_208_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_208_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_208_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_208_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_208_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_208_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_208_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_208_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_208_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_208_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_208_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_208_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_208_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_208_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_208_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_208_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_208_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_208_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_208_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_208_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_208_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_208_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_208_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_208_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_208_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_208_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_209 ( // @[mac.scala 29:63]
    .clock(PECross_209_clock),
    .reset(PECross_209_reset),
    .multiply_io_input_io_sumIn_ready(PECross_209_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_209_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_209_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_209_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_209_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_209_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_209_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_209_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_209_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_209_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_209_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_209_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_209_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_209_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_209_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_209_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_209_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_209_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_209_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_209_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_209_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_209_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_209_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_209_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_209_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_209_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_209_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_210 ( // @[mac.scala 29:63]
    .clock(PECross_210_clock),
    .reset(PECross_210_reset),
    .multiply_io_input_io_sumIn_ready(PECross_210_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_210_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_210_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_210_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_210_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_210_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_210_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_210_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_210_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_210_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_210_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_210_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_210_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_210_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_210_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_210_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_210_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_210_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_210_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_210_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_210_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_210_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_210_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_210_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_210_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_210_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_210_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_211 ( // @[mac.scala 29:63]
    .clock(PECross_211_clock),
    .reset(PECross_211_reset),
    .multiply_io_input_io_sumIn_ready(PECross_211_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_211_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_211_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_211_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_211_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_211_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_211_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_211_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_211_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_211_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_211_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_211_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_211_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_211_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_211_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_211_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_211_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_211_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_211_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_211_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_211_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_211_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_211_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_211_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_211_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_211_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_211_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_212 ( // @[mac.scala 29:63]
    .clock(PECross_212_clock),
    .reset(PECross_212_reset),
    .multiply_io_input_io_sumIn_ready(PECross_212_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_212_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_212_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_212_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_212_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_212_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_212_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_212_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_212_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_212_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_212_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_212_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_212_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_212_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_212_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_212_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_212_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_212_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_212_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_212_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_212_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_212_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_212_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_212_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_212_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_212_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_212_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_213 ( // @[mac.scala 29:63]
    .clock(PECross_213_clock),
    .reset(PECross_213_reset),
    .multiply_io_input_io_sumIn_ready(PECross_213_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_213_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_213_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_213_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_213_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_213_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_213_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_213_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_213_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_213_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_213_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_213_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_213_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_213_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_213_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_213_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_213_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_213_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_213_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_213_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_213_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_213_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_213_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_213_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_213_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_213_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_213_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_214 ( // @[mac.scala 29:63]
    .clock(PECross_214_clock),
    .reset(PECross_214_reset),
    .multiply_io_input_io_sumIn_ready(PECross_214_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_214_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_214_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_214_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_214_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_214_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_214_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_214_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_214_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_214_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_214_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_214_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_214_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_214_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_214_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_214_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_214_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_214_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_214_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_214_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_214_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_214_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_214_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_214_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_214_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_214_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_214_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_215 ( // @[mac.scala 29:63]
    .clock(PECross_215_clock),
    .reset(PECross_215_reset),
    .multiply_io_input_io_sumIn_ready(PECross_215_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_215_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_215_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_215_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_215_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_215_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_215_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_215_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_215_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_215_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_215_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_215_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_215_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_215_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_215_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_215_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_215_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_215_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_215_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_215_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_215_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_215_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_215_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_215_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_215_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_215_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_215_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_216 ( // @[mac.scala 29:63]
    .clock(PECross_216_clock),
    .reset(PECross_216_reset),
    .multiply_io_input_io_sumIn_ready(PECross_216_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_216_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_216_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_216_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_216_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_216_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_216_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_216_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_216_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_216_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_216_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_216_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_216_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_216_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_216_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_216_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_216_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_216_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_216_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_216_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_216_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_216_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_216_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_216_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_216_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_216_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_216_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_217 ( // @[mac.scala 29:63]
    .clock(PECross_217_clock),
    .reset(PECross_217_reset),
    .multiply_io_input_io_sumIn_ready(PECross_217_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_217_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_217_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_217_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_217_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_217_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_217_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_217_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_217_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_217_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_217_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_217_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_217_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_217_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_217_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_217_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_217_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_217_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_217_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_217_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_217_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_217_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_217_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_217_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_217_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_217_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_217_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_218 ( // @[mac.scala 29:63]
    .clock(PECross_218_clock),
    .reset(PECross_218_reset),
    .multiply_io_input_io_sumIn_ready(PECross_218_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_218_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_218_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_218_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_218_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_218_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_218_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_218_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_218_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_218_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_218_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_218_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_218_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_218_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_218_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_218_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_218_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_218_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_218_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_218_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_218_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_218_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_218_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_218_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_218_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_218_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_218_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_219 ( // @[mac.scala 29:63]
    .clock(PECross_219_clock),
    .reset(PECross_219_reset),
    .multiply_io_input_io_sumIn_ready(PECross_219_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_219_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_219_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_219_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_219_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_219_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_219_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_219_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_219_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_219_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_219_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_219_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_219_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_219_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_219_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_219_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_219_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_219_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_219_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_219_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_219_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_219_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_219_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_219_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_219_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_219_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_219_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_220 ( // @[mac.scala 29:63]
    .clock(PECross_220_clock),
    .reset(PECross_220_reset),
    .multiply_io_input_io_sumIn_ready(PECross_220_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_220_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_220_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_220_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_220_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_220_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_220_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_220_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_220_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_220_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_220_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_220_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_220_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_220_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_220_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_220_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_220_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_220_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_220_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_220_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_220_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_220_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_220_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_220_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_220_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_220_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_220_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_221 ( // @[mac.scala 29:63]
    .clock(PECross_221_clock),
    .reset(PECross_221_reset),
    .multiply_io_input_io_sumIn_ready(PECross_221_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_221_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_221_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_221_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_221_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_221_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_221_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_221_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_221_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_221_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_221_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_221_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_221_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_221_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_221_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_221_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_221_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_221_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_221_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_221_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_221_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_221_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_221_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_221_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_221_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_221_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_221_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_222 ( // @[mac.scala 29:63]
    .clock(PECross_222_clock),
    .reset(PECross_222_reset),
    .multiply_io_input_io_sumIn_ready(PECross_222_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_222_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_222_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_222_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_222_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_222_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_222_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_222_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_222_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_222_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_222_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_222_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_222_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_222_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_222_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_222_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_222_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_222_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_222_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_222_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_222_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_222_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_222_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_222_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_222_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_222_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_222_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_223 ( // @[mac.scala 29:63]
    .clock(PECross_223_clock),
    .reset(PECross_223_reset),
    .multiply_io_input_io_sumIn_ready(PECross_223_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_223_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_223_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_223_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_223_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_223_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_223_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_223_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_223_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_223_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_223_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_223_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_223_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_223_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_223_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_223_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_223_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_223_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_223_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_223_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_223_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_223_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_223_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_223_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_223_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_223_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_223_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_224 ( // @[mac.scala 29:63]
    .clock(PECross_224_clock),
    .reset(PECross_224_reset),
    .multiply_io_input_io_sumIn_ready(PECross_224_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_224_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_224_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_224_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_224_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_224_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_224_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_224_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_224_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_224_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_224_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_224_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_224_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_224_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_224_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_224_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_224_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_224_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_224_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_224_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_224_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_224_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_224_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_224_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_224_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_224_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_224_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_225 ( // @[mac.scala 29:63]
    .clock(PECross_225_clock),
    .reset(PECross_225_reset),
    .multiply_io_input_io_sumIn_ready(PECross_225_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_225_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_225_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_225_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_225_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_225_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_225_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_225_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_225_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_225_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_225_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_225_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_225_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_225_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_225_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_225_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_225_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_225_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_225_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_225_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_225_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_225_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_225_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_225_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_225_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_225_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_225_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_226 ( // @[mac.scala 29:63]
    .clock(PECross_226_clock),
    .reset(PECross_226_reset),
    .multiply_io_input_io_sumIn_ready(PECross_226_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_226_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_226_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_226_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_226_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_226_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_226_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_226_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_226_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_226_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_226_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_226_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_226_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_226_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_226_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_226_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_226_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_226_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_226_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_226_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_226_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_226_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_226_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_226_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_226_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_226_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_226_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_227 ( // @[mac.scala 29:63]
    .clock(PECross_227_clock),
    .reset(PECross_227_reset),
    .multiply_io_input_io_sumIn_ready(PECross_227_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_227_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_227_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_227_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_227_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_227_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_227_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_227_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_227_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_227_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_227_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_227_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_227_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_227_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_227_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_227_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_227_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_227_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_227_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_227_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_227_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_227_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_227_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_227_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_227_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_227_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_227_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_228 ( // @[mac.scala 29:63]
    .clock(PECross_228_clock),
    .reset(PECross_228_reset),
    .multiply_io_input_io_sumIn_ready(PECross_228_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_228_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_228_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_228_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_228_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_228_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_228_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_228_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_228_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_228_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_228_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_228_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_228_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_228_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_228_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_228_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_228_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_228_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_228_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_228_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_228_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_228_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_228_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_228_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_228_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_228_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_228_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_229 ( // @[mac.scala 29:63]
    .clock(PECross_229_clock),
    .reset(PECross_229_reset),
    .multiply_io_input_io_sumIn_ready(PECross_229_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_229_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_229_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_229_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_229_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_229_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_229_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_229_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_229_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_229_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_229_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_229_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_229_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_229_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_229_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_229_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_229_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_229_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_229_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_229_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_229_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_229_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_229_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_229_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_229_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_229_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_229_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_230 ( // @[mac.scala 29:63]
    .clock(PECross_230_clock),
    .reset(PECross_230_reset),
    .multiply_io_input_io_sumIn_ready(PECross_230_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_230_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_230_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_230_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_230_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_230_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_230_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_230_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_230_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_230_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_230_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_230_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_230_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_230_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_230_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_230_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_230_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_230_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_230_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_230_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_230_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_230_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_230_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_230_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_230_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_230_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_230_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_231 ( // @[mac.scala 29:63]
    .clock(PECross_231_clock),
    .reset(PECross_231_reset),
    .multiply_io_input_io_sumIn_ready(PECross_231_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_231_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_231_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_231_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_231_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_231_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_231_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_231_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_231_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_231_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_231_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_231_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_231_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_231_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_231_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_231_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_231_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_231_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_231_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_231_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_231_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_231_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_231_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_231_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_231_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_231_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_231_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_232 ( // @[mac.scala 29:63]
    .clock(PECross_232_clock),
    .reset(PECross_232_reset),
    .multiply_io_input_io_sumIn_ready(PECross_232_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_232_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_232_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_232_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_232_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_232_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_232_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_232_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_232_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_232_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_232_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_232_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_232_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_232_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_232_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_232_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_232_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_232_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_232_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_232_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_232_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_232_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_232_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_232_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_232_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_232_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_232_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_233 ( // @[mac.scala 29:63]
    .clock(PECross_233_clock),
    .reset(PECross_233_reset),
    .multiply_io_input_io_sumIn_ready(PECross_233_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_233_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_233_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_233_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_233_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_233_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_233_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_233_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_233_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_233_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_233_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_233_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_233_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_233_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_233_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_233_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_233_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_233_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_233_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_233_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_233_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_233_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_233_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_233_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_233_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_233_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_233_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_234 ( // @[mac.scala 29:63]
    .clock(PECross_234_clock),
    .reset(PECross_234_reset),
    .multiply_io_input_io_sumIn_ready(PECross_234_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_234_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_234_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_234_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_234_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_234_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_234_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_234_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_234_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_234_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_234_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_234_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_234_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_234_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_234_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_234_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_234_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_234_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_234_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_234_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_234_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_234_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_234_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_234_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_234_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_234_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_234_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_235 ( // @[mac.scala 29:63]
    .clock(PECross_235_clock),
    .reset(PECross_235_reset),
    .multiply_io_input_io_sumIn_ready(PECross_235_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_235_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_235_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_235_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_235_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_235_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_235_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_235_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_235_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_235_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_235_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_235_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_235_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_235_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_235_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_235_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_235_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_235_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_235_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_235_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_235_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_235_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_235_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_235_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_235_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_235_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_235_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_236 ( // @[mac.scala 29:63]
    .clock(PECross_236_clock),
    .reset(PECross_236_reset),
    .multiply_io_input_io_sumIn_ready(PECross_236_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_236_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_236_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_236_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_236_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_236_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_236_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_236_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_236_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_236_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_236_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_236_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_236_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_236_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_236_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_236_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_236_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_236_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_236_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_236_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_236_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_236_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_236_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_236_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_236_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_236_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_236_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_237 ( // @[mac.scala 29:63]
    .clock(PECross_237_clock),
    .reset(PECross_237_reset),
    .multiply_io_input_io_sumIn_ready(PECross_237_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_237_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_237_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_237_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_237_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_237_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_237_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_237_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_237_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_237_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_237_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_237_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_237_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_237_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_237_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_237_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_237_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_237_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_237_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_237_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_237_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_237_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_237_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_237_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_237_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_237_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_237_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_238 ( // @[mac.scala 29:63]
    .clock(PECross_238_clock),
    .reset(PECross_238_reset),
    .multiply_io_input_io_sumIn_ready(PECross_238_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_238_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_238_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_238_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_238_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_238_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_238_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_238_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_238_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_238_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_238_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_238_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_238_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_238_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_238_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_238_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_238_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_238_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_238_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_238_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_238_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_238_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_238_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_238_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_238_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_238_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_238_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_239 ( // @[mac.scala 29:63]
    .clock(PECross_239_clock),
    .reset(PECross_239_reset),
    .multiply_io_input_io_sumIn_ready(PECross_239_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_239_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_239_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_239_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_239_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_239_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_239_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_239_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_239_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_239_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_239_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_239_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_239_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_239_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_239_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_239_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_239_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_239_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_239_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_239_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_239_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_239_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_239_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_239_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_239_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_239_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_239_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_240 ( // @[mac.scala 29:63]
    .clock(PECross_240_clock),
    .reset(PECross_240_reset),
    .multiply_io_input_io_sumIn_ready(PECross_240_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_240_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_240_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_240_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_240_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_240_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_240_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_240_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_240_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_240_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_240_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_240_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_240_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_240_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_240_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_240_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_240_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_240_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_240_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_240_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_240_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_240_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_240_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_240_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_240_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_240_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_240_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_241 ( // @[mac.scala 29:63]
    .clock(PECross_241_clock),
    .reset(PECross_241_reset),
    .multiply_io_input_io_sumIn_ready(PECross_241_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_241_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_241_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_241_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_241_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_241_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_241_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_241_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_241_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_241_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_241_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_241_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_241_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_241_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_241_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_241_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_241_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_241_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_241_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_241_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_241_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_241_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_241_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_241_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_241_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_241_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_241_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_242 ( // @[mac.scala 29:63]
    .clock(PECross_242_clock),
    .reset(PECross_242_reset),
    .multiply_io_input_io_sumIn_ready(PECross_242_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_242_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_242_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_242_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_242_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_242_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_242_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_242_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_242_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_242_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_242_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_242_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_242_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_242_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_242_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_242_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_242_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_242_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_242_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_242_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_242_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_242_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_242_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_242_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_242_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_242_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_242_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_243 ( // @[mac.scala 29:63]
    .clock(PECross_243_clock),
    .reset(PECross_243_reset),
    .multiply_io_input_io_sumIn_ready(PECross_243_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_243_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_243_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_243_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_243_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_243_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_243_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_243_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_243_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_243_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_243_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_243_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_243_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_243_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_243_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_243_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_243_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_243_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_243_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_243_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_243_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_243_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_243_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_243_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_243_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_243_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_243_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_244 ( // @[mac.scala 29:63]
    .clock(PECross_244_clock),
    .reset(PECross_244_reset),
    .multiply_io_input_io_sumIn_ready(PECross_244_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_244_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_244_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_244_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_244_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_244_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_244_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_244_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_244_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_244_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_244_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_244_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_244_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_244_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_244_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_244_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_244_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_244_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_244_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_244_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_244_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_244_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_244_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_244_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_244_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_244_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_244_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_245 ( // @[mac.scala 29:63]
    .clock(PECross_245_clock),
    .reset(PECross_245_reset),
    .multiply_io_input_io_sumIn_ready(PECross_245_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_245_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_245_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_245_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_245_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_245_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_245_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_245_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_245_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_245_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_245_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_245_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_245_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_245_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_245_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_245_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_245_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_245_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_245_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_245_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_245_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_245_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_245_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_245_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_245_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_245_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_245_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_246 ( // @[mac.scala 29:63]
    .clock(PECross_246_clock),
    .reset(PECross_246_reset),
    .multiply_io_input_io_sumIn_ready(PECross_246_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_246_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_246_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_246_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_246_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_246_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_246_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_246_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_246_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_246_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_246_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_246_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_246_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_246_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_246_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_246_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_246_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_246_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_246_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_246_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_246_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_246_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_246_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_246_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_246_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_246_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_246_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_247 ( // @[mac.scala 29:63]
    .clock(PECross_247_clock),
    .reset(PECross_247_reset),
    .multiply_io_input_io_sumIn_ready(PECross_247_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_247_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_247_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_247_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_247_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_247_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_247_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_247_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_247_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_247_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_247_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_247_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_247_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_247_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_247_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_247_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_247_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_247_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_247_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_247_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_247_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_247_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_247_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_247_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_247_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_247_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_247_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_248 ( // @[mac.scala 29:63]
    .clock(PECross_248_clock),
    .reset(PECross_248_reset),
    .multiply_io_input_io_sumIn_ready(PECross_248_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_248_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_248_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_248_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_248_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_248_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_248_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_248_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_248_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_248_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_248_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_248_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_248_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_248_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_248_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_248_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_248_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_248_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_248_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_248_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_248_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_248_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_248_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_248_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_248_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_248_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_248_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_249 ( // @[mac.scala 29:63]
    .clock(PECross_249_clock),
    .reset(PECross_249_reset),
    .multiply_io_input_io_sumIn_ready(PECross_249_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_249_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_249_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_249_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_249_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_249_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_249_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_249_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_249_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_249_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_249_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_249_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_249_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_249_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_249_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_249_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_249_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_249_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_249_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_249_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_249_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_249_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_249_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_249_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_249_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_249_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_249_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_250 ( // @[mac.scala 29:63]
    .clock(PECross_250_clock),
    .reset(PECross_250_reset),
    .multiply_io_input_io_sumIn_ready(PECross_250_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_250_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_250_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_250_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_250_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_250_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_250_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_250_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_250_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_250_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_250_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_250_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_250_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_250_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_250_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_250_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_250_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_250_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_250_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_250_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_250_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_250_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_250_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_250_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_250_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_250_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_250_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_251 ( // @[mac.scala 29:63]
    .clock(PECross_251_clock),
    .reset(PECross_251_reset),
    .multiply_io_input_io_sumIn_ready(PECross_251_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_251_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_251_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_251_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_251_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_251_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_251_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_251_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_251_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_251_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_251_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_251_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_251_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_251_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_251_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_251_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_251_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_251_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_251_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_251_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_251_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_251_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_251_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_251_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_251_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_251_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_251_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_252 ( // @[mac.scala 29:63]
    .clock(PECross_252_clock),
    .reset(PECross_252_reset),
    .multiply_io_input_io_sumIn_ready(PECross_252_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_252_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_252_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_252_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_252_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_252_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_252_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_252_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_252_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_252_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_252_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_252_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_252_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_252_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_252_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_252_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_252_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_252_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_252_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_252_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_252_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_252_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_252_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_252_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_252_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_252_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_252_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_253 ( // @[mac.scala 29:63]
    .clock(PECross_253_clock),
    .reset(PECross_253_reset),
    .multiply_io_input_io_sumIn_ready(PECross_253_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_253_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_253_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_253_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_253_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_253_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_253_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_253_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_253_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_253_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_253_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_253_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_253_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_253_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_253_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_253_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_253_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_253_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_253_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_253_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_253_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_253_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_253_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_253_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_253_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_253_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_253_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_254 ( // @[mac.scala 29:63]
    .clock(PECross_254_clock),
    .reset(PECross_254_reset),
    .multiply_io_input_io_sumIn_ready(PECross_254_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_254_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_254_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_254_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_254_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_254_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_254_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_254_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_254_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_254_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_254_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_254_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_254_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_254_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_254_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_254_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_254_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_254_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_254_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_254_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_254_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_254_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_254_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_254_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_254_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_254_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_254_multiply_io_input_io_weiOut_bits_last)
  );
  PECross PECross_255 ( // @[mac.scala 29:63]
    .clock(PECross_255_clock),
    .reset(PECross_255_reset),
    .multiply_io_input_io_sumIn_ready(PECross_255_multiply_io_input_io_sumIn_ready),
    .multiply_io_input_io_sumIn_valid(PECross_255_multiply_io_input_io_sumIn_valid),
    .multiply_io_input_io_sumIn_bits_x_0(PECross_255_multiply_io_input_io_sumIn_bits_x_0),
    .multiply_io_input_io_sumIn_bits_last(PECross_255_multiply_io_input_io_sumIn_bits_last),
    .multiply_io_input_io_sumOut_ready(PECross_255_multiply_io_input_io_sumOut_ready),
    .multiply_io_input_io_sumOut_valid(PECross_255_multiply_io_input_io_sumOut_valid),
    .multiply_io_input_io_sumOut_bits_x_0(PECross_255_multiply_io_input_io_sumOut_bits_x_0),
    .multiply_io_input_io_sumOut_bits_last(PECross_255_multiply_io_input_io_sumOut_bits_last),
    .multiply_io_input_io_statSel(PECross_255_multiply_io_input_io_statSel),
    .multiply_io_input_io_weiEn(PECross_255_multiply_io_input_io_weiEn),
    .multiply_io_input_io_actEn(PECross_255_multiply_io_input_io_actEn),
    .multiply_io_input_io_actIn_ready(PECross_255_multiply_io_input_io_actIn_ready),
    .multiply_io_input_io_actIn_valid(PECross_255_multiply_io_input_io_actIn_valid),
    .multiply_io_input_io_actIn_bits_x_0(PECross_255_multiply_io_input_io_actIn_bits_x_0),
    .multiply_io_input_io_actIn_bits_last(PECross_255_multiply_io_input_io_actIn_bits_last),
    .multiply_io_input_io_weiIn_ready(PECross_255_multiply_io_input_io_weiIn_ready),
    .multiply_io_input_io_weiIn_valid(PECross_255_multiply_io_input_io_weiIn_valid),
    .multiply_io_input_io_weiIn_bits_x_0(PECross_255_multiply_io_input_io_weiIn_bits_x_0),
    .multiply_io_input_io_weiIn_bits_last(PECross_255_multiply_io_input_io_weiIn_bits_last),
    .multiply_io_input_io_actOut_ready(PECross_255_multiply_io_input_io_actOut_ready),
    .multiply_io_input_io_actOut_valid(PECross_255_multiply_io_input_io_actOut_valid),
    .multiply_io_input_io_actOut_bits_x_0(PECross_255_multiply_io_input_io_actOut_bits_x_0),
    .multiply_io_input_io_actOut_bits_last(PECross_255_multiply_io_input_io_actOut_bits_last),
    .multiply_io_input_io_weiOut_ready(PECross_255_multiply_io_input_io_weiOut_ready),
    .multiply_io_input_io_weiOut_valid(PECross_255_multiply_io_input_io_weiOut_valid),
    .multiply_io_input_io_weiOut_bits_x_0(PECross_255_multiply_io_input_io_weiOut_bits_x_0),
    .multiply_io_input_io_weiOut_bits_last(PECross_255_multiply_io_input_io_weiOut_bits_last)
  );
  assign io_actIn_0_ready = PECross_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_1_ready = PECross_16_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_2_ready = PECross_32_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_3_ready = PECross_48_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_4_ready = PECross_64_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_5_ready = PECross_80_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_6_ready = PECross_96_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_7_ready = PECross_112_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_8_ready = PECross_128_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_9_ready = PECross_144_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_10_ready = PECross_160_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_11_ready = PECross_176_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_12_ready = PECross_192_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_13_ready = PECross_208_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_14_ready = PECross_224_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_actIn_15_ready = PECross_240_multiply_io_input_io_actIn_ready; // @[mac.scala 32:28]
  assign io_weiIn_0_ready = PECross_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_1_ready = PECross_1_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_2_ready = PECross_2_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_3_ready = PECross_3_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_4_ready = PECross_4_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_5_ready = PECross_5_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_6_ready = PECross_6_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_7_ready = PECross_7_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_8_ready = PECross_8_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_9_ready = PECross_9_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_10_ready = PECross_10_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_11_ready = PECross_11_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_12_ready = PECross_12_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_13_ready = PECross_13_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_14_ready = PECross_14_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_weiIn_15_ready = PECross_15_multiply_io_input_io_weiIn_ready; // @[mac.scala 40:28]
  assign io_sumIn_0_ready = PECross_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_1_ready = PECross_16_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_2_ready = PECross_32_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_3_ready = PECross_48_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_4_ready = PECross_64_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_5_ready = PECross_80_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_6_ready = PECross_96_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_7_ready = PECross_112_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_8_ready = PECross_128_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_9_ready = PECross_144_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_10_ready = PECross_160_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_11_ready = PECross_176_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_12_ready = PECross_192_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_13_ready = PECross_208_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_14_ready = PECross_224_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumIn_15_ready = PECross_240_multiply_io_input_io_sumIn_ready; // @[mac.scala 33:28]
  assign io_sumOut_0_valid = PECross_15_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_0_bits_x_0 = PECross_15_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_0_bits_last = PECross_15_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_1_valid = PECross_31_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_1_bits_x_0 = PECross_31_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_1_bits_last = PECross_31_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_2_valid = PECross_47_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_2_bits_x_0 = PECross_47_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_2_bits_last = PECross_47_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_3_valid = PECross_63_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_3_bits_x_0 = PECross_63_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_3_bits_last = PECross_63_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_4_valid = PECross_79_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_4_bits_x_0 = PECross_79_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_4_bits_last = PECross_79_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_5_valid = PECross_95_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_5_bits_x_0 = PECross_95_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_5_bits_last = PECross_95_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_6_valid = PECross_111_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_6_bits_x_0 = PECross_111_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_6_bits_last = PECross_111_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_7_valid = PECross_127_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_7_bits_x_0 = PECross_127_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_7_bits_last = PECross_127_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_8_valid = PECross_143_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_8_bits_x_0 = PECross_143_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_8_bits_last = PECross_143_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_9_valid = PECross_159_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_9_bits_x_0 = PECross_159_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_9_bits_last = PECross_159_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_10_valid = PECross_175_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_10_bits_x_0 = PECross_175_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_10_bits_last = PECross_175_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_11_valid = PECross_191_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_11_bits_x_0 = PECross_191_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_11_bits_last = PECross_191_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_12_valid = PECross_207_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_12_bits_x_0 = PECross_207_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_12_bits_last = PECross_207_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_13_valid = PECross_223_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_13_bits_x_0 = PECross_223_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_13_bits_last = PECross_223_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_14_valid = PECross_239_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_14_bits_x_0 = PECross_239_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_14_bits_last = PECross_239_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign io_sumOut_15_valid = PECross_255_multiply_io_input_io_sumOut_valid; // @[mac.scala 45:29]
  assign io_sumOut_15_bits_x_0 = PECross_255_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 45:29]
  assign io_sumOut_15_bits_last = PECross_255_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 45:29]
  assign PECross_clock = clock;
  assign PECross_reset = rst;
  assign PECross_multiply_io_input_io_sumIn_valid = io_sumIn_0_valid; // @[mac.scala 33:28]
  assign PECross_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_0_bits_x_0; // @[mac.scala 33:28]
  assign PECross_multiply_io_input_io_sumIn_bits_last = io_sumIn_0_bits_last; // @[mac.scala 33:28]
  assign PECross_multiply_io_input_io_sumOut_ready = PECross_1_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_multiply_io_input_io_actIn_valid = io_actIn_0_valid; // @[mac.scala 32:28]
  assign PECross_multiply_io_input_io_actIn_bits_x_0 = io_actIn_0_bits_x_0; // @[mac.scala 32:28]
  assign PECross_multiply_io_input_io_actIn_bits_last = io_actIn_0_bits_last; // @[mac.scala 32:28]
  assign PECross_multiply_io_input_io_weiIn_valid = io_weiIn_0_valid; // @[mac.scala 40:28]
  assign PECross_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_0_bits_x_0; // @[mac.scala 40:28]
  assign PECross_multiply_io_input_io_weiIn_bits_last = io_weiIn_0_bits_last; // @[mac.scala 40:28]
  assign PECross_multiply_io_input_io_actOut_ready = PECross_1_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_multiply_io_input_io_weiOut_ready = PECross_16_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_1_clock = clock;
  assign PECross_1_reset = rst;
  assign PECross_1_multiply_io_input_io_sumIn_valid = PECross_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_1_multiply_io_input_io_sumIn_bits_x_0 = PECross_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_1_multiply_io_input_io_sumIn_bits_last = PECross_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_1_multiply_io_input_io_sumOut_ready = PECross_2_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_1_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_1_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_1_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_1_multiply_io_input_io_actIn_valid = PECross_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_1_multiply_io_input_io_actIn_bits_x_0 = PECross_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_1_multiply_io_input_io_actIn_bits_last = PECross_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_1_multiply_io_input_io_weiIn_valid = io_weiIn_1_valid; // @[mac.scala 40:28]
  assign PECross_1_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_1_bits_x_0; // @[mac.scala 40:28]
  assign PECross_1_multiply_io_input_io_weiIn_bits_last = io_weiIn_1_bits_last; // @[mac.scala 40:28]
  assign PECross_1_multiply_io_input_io_actOut_ready = PECross_2_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_1_multiply_io_input_io_weiOut_ready = PECross_17_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_2_clock = clock;
  assign PECross_2_reset = rst;
  assign PECross_2_multiply_io_input_io_sumIn_valid = PECross_1_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_2_multiply_io_input_io_sumIn_bits_x_0 = PECross_1_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_2_multiply_io_input_io_sumIn_bits_last = PECross_1_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_2_multiply_io_input_io_sumOut_ready = PECross_3_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_2_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_2_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_2_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_2_multiply_io_input_io_actIn_valid = PECross_1_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_2_multiply_io_input_io_actIn_bits_x_0 = PECross_1_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_2_multiply_io_input_io_actIn_bits_last = PECross_1_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_2_multiply_io_input_io_weiIn_valid = io_weiIn_2_valid; // @[mac.scala 40:28]
  assign PECross_2_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_2_bits_x_0; // @[mac.scala 40:28]
  assign PECross_2_multiply_io_input_io_weiIn_bits_last = io_weiIn_2_bits_last; // @[mac.scala 40:28]
  assign PECross_2_multiply_io_input_io_actOut_ready = PECross_3_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_2_multiply_io_input_io_weiOut_ready = PECross_18_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_3_clock = clock;
  assign PECross_3_reset = rst;
  assign PECross_3_multiply_io_input_io_sumIn_valid = PECross_2_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_3_multiply_io_input_io_sumIn_bits_x_0 = PECross_2_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_3_multiply_io_input_io_sumIn_bits_last = PECross_2_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_3_multiply_io_input_io_sumOut_ready = PECross_4_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_3_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_3_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_3_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_3_multiply_io_input_io_actIn_valid = PECross_2_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_3_multiply_io_input_io_actIn_bits_x_0 = PECross_2_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_3_multiply_io_input_io_actIn_bits_last = PECross_2_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_3_multiply_io_input_io_weiIn_valid = io_weiIn_3_valid; // @[mac.scala 40:28]
  assign PECross_3_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_3_bits_x_0; // @[mac.scala 40:28]
  assign PECross_3_multiply_io_input_io_weiIn_bits_last = io_weiIn_3_bits_last; // @[mac.scala 40:28]
  assign PECross_3_multiply_io_input_io_actOut_ready = PECross_4_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_3_multiply_io_input_io_weiOut_ready = PECross_19_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_4_clock = clock;
  assign PECross_4_reset = rst;
  assign PECross_4_multiply_io_input_io_sumIn_valid = PECross_3_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_4_multiply_io_input_io_sumIn_bits_x_0 = PECross_3_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_4_multiply_io_input_io_sumIn_bits_last = PECross_3_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_4_multiply_io_input_io_sumOut_ready = PECross_5_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_4_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_4_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_4_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_4_multiply_io_input_io_actIn_valid = PECross_3_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_4_multiply_io_input_io_actIn_bits_x_0 = PECross_3_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_4_multiply_io_input_io_actIn_bits_last = PECross_3_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_4_multiply_io_input_io_weiIn_valid = io_weiIn_4_valid; // @[mac.scala 40:28]
  assign PECross_4_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_4_bits_x_0; // @[mac.scala 40:28]
  assign PECross_4_multiply_io_input_io_weiIn_bits_last = io_weiIn_4_bits_last; // @[mac.scala 40:28]
  assign PECross_4_multiply_io_input_io_actOut_ready = PECross_5_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_4_multiply_io_input_io_weiOut_ready = PECross_20_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_5_clock = clock;
  assign PECross_5_reset = rst;
  assign PECross_5_multiply_io_input_io_sumIn_valid = PECross_4_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_5_multiply_io_input_io_sumIn_bits_x_0 = PECross_4_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_5_multiply_io_input_io_sumIn_bits_last = PECross_4_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_5_multiply_io_input_io_sumOut_ready = PECross_6_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_5_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_5_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_5_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_5_multiply_io_input_io_actIn_valid = PECross_4_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_5_multiply_io_input_io_actIn_bits_x_0 = PECross_4_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_5_multiply_io_input_io_actIn_bits_last = PECross_4_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_5_multiply_io_input_io_weiIn_valid = io_weiIn_5_valid; // @[mac.scala 40:28]
  assign PECross_5_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_5_bits_x_0; // @[mac.scala 40:28]
  assign PECross_5_multiply_io_input_io_weiIn_bits_last = io_weiIn_5_bits_last; // @[mac.scala 40:28]
  assign PECross_5_multiply_io_input_io_actOut_ready = PECross_6_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_5_multiply_io_input_io_weiOut_ready = PECross_21_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_6_clock = clock;
  assign PECross_6_reset = rst;
  assign PECross_6_multiply_io_input_io_sumIn_valid = PECross_5_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_6_multiply_io_input_io_sumIn_bits_x_0 = PECross_5_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_6_multiply_io_input_io_sumIn_bits_last = PECross_5_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_6_multiply_io_input_io_sumOut_ready = PECross_7_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_6_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_6_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_6_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_6_multiply_io_input_io_actIn_valid = PECross_5_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_6_multiply_io_input_io_actIn_bits_x_0 = PECross_5_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_6_multiply_io_input_io_actIn_bits_last = PECross_5_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_6_multiply_io_input_io_weiIn_valid = io_weiIn_6_valid; // @[mac.scala 40:28]
  assign PECross_6_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_6_bits_x_0; // @[mac.scala 40:28]
  assign PECross_6_multiply_io_input_io_weiIn_bits_last = io_weiIn_6_bits_last; // @[mac.scala 40:28]
  assign PECross_6_multiply_io_input_io_actOut_ready = PECross_7_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_6_multiply_io_input_io_weiOut_ready = PECross_22_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_7_clock = clock;
  assign PECross_7_reset = rst;
  assign PECross_7_multiply_io_input_io_sumIn_valid = PECross_6_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_7_multiply_io_input_io_sumIn_bits_x_0 = PECross_6_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_7_multiply_io_input_io_sumIn_bits_last = PECross_6_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_7_multiply_io_input_io_sumOut_ready = PECross_8_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_7_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_7_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_7_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_7_multiply_io_input_io_actIn_valid = PECross_6_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_7_multiply_io_input_io_actIn_bits_x_0 = PECross_6_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_7_multiply_io_input_io_actIn_bits_last = PECross_6_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_7_multiply_io_input_io_weiIn_valid = io_weiIn_7_valid; // @[mac.scala 40:28]
  assign PECross_7_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_7_bits_x_0; // @[mac.scala 40:28]
  assign PECross_7_multiply_io_input_io_weiIn_bits_last = io_weiIn_7_bits_last; // @[mac.scala 40:28]
  assign PECross_7_multiply_io_input_io_actOut_ready = PECross_8_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_7_multiply_io_input_io_weiOut_ready = PECross_23_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_8_clock = clock;
  assign PECross_8_reset = rst;
  assign PECross_8_multiply_io_input_io_sumIn_valid = PECross_7_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_8_multiply_io_input_io_sumIn_bits_x_0 = PECross_7_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_8_multiply_io_input_io_sumIn_bits_last = PECross_7_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_8_multiply_io_input_io_sumOut_ready = PECross_9_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_8_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_8_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_8_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_8_multiply_io_input_io_actIn_valid = PECross_7_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_8_multiply_io_input_io_actIn_bits_x_0 = PECross_7_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_8_multiply_io_input_io_actIn_bits_last = PECross_7_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_8_multiply_io_input_io_weiIn_valid = io_weiIn_8_valid; // @[mac.scala 40:28]
  assign PECross_8_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_8_bits_x_0; // @[mac.scala 40:28]
  assign PECross_8_multiply_io_input_io_weiIn_bits_last = io_weiIn_8_bits_last; // @[mac.scala 40:28]
  assign PECross_8_multiply_io_input_io_actOut_ready = PECross_9_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_8_multiply_io_input_io_weiOut_ready = PECross_24_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_9_clock = clock;
  assign PECross_9_reset = rst;
  assign PECross_9_multiply_io_input_io_sumIn_valid = PECross_8_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_9_multiply_io_input_io_sumIn_bits_x_0 = PECross_8_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_9_multiply_io_input_io_sumIn_bits_last = PECross_8_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_9_multiply_io_input_io_sumOut_ready = PECross_10_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_9_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_9_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_9_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_9_multiply_io_input_io_actIn_valid = PECross_8_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_9_multiply_io_input_io_actIn_bits_x_0 = PECross_8_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_9_multiply_io_input_io_actIn_bits_last = PECross_8_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_9_multiply_io_input_io_weiIn_valid = io_weiIn_9_valid; // @[mac.scala 40:28]
  assign PECross_9_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_9_bits_x_0; // @[mac.scala 40:28]
  assign PECross_9_multiply_io_input_io_weiIn_bits_last = io_weiIn_9_bits_last; // @[mac.scala 40:28]
  assign PECross_9_multiply_io_input_io_actOut_ready = PECross_10_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_9_multiply_io_input_io_weiOut_ready = PECross_25_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_10_clock = clock;
  assign PECross_10_reset = rst;
  assign PECross_10_multiply_io_input_io_sumIn_valid = PECross_9_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_10_multiply_io_input_io_sumIn_bits_x_0 = PECross_9_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_10_multiply_io_input_io_sumIn_bits_last = PECross_9_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_10_multiply_io_input_io_sumOut_ready = PECross_11_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_10_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_10_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_10_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_10_multiply_io_input_io_actIn_valid = PECross_9_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_10_multiply_io_input_io_actIn_bits_x_0 = PECross_9_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_10_multiply_io_input_io_actIn_bits_last = PECross_9_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_10_multiply_io_input_io_weiIn_valid = io_weiIn_10_valid; // @[mac.scala 40:28]
  assign PECross_10_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_10_bits_x_0; // @[mac.scala 40:28]
  assign PECross_10_multiply_io_input_io_weiIn_bits_last = io_weiIn_10_bits_last; // @[mac.scala 40:28]
  assign PECross_10_multiply_io_input_io_actOut_ready = PECross_11_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_10_multiply_io_input_io_weiOut_ready = PECross_26_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_11_clock = clock;
  assign PECross_11_reset = rst;
  assign PECross_11_multiply_io_input_io_sumIn_valid = PECross_10_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_11_multiply_io_input_io_sumIn_bits_x_0 = PECross_10_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_11_multiply_io_input_io_sumIn_bits_last = PECross_10_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_11_multiply_io_input_io_sumOut_ready = PECross_12_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_11_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_11_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_11_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_11_multiply_io_input_io_actIn_valid = PECross_10_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_11_multiply_io_input_io_actIn_bits_x_0 = PECross_10_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_11_multiply_io_input_io_actIn_bits_last = PECross_10_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_11_multiply_io_input_io_weiIn_valid = io_weiIn_11_valid; // @[mac.scala 40:28]
  assign PECross_11_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_11_bits_x_0; // @[mac.scala 40:28]
  assign PECross_11_multiply_io_input_io_weiIn_bits_last = io_weiIn_11_bits_last; // @[mac.scala 40:28]
  assign PECross_11_multiply_io_input_io_actOut_ready = PECross_12_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_11_multiply_io_input_io_weiOut_ready = PECross_27_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_12_clock = clock;
  assign PECross_12_reset = rst;
  assign PECross_12_multiply_io_input_io_sumIn_valid = PECross_11_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_12_multiply_io_input_io_sumIn_bits_x_0 = PECross_11_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_12_multiply_io_input_io_sumIn_bits_last = PECross_11_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_12_multiply_io_input_io_sumOut_ready = PECross_13_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_12_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_12_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_12_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_12_multiply_io_input_io_actIn_valid = PECross_11_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_12_multiply_io_input_io_actIn_bits_x_0 = PECross_11_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_12_multiply_io_input_io_actIn_bits_last = PECross_11_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_12_multiply_io_input_io_weiIn_valid = io_weiIn_12_valid; // @[mac.scala 40:28]
  assign PECross_12_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_12_bits_x_0; // @[mac.scala 40:28]
  assign PECross_12_multiply_io_input_io_weiIn_bits_last = io_weiIn_12_bits_last; // @[mac.scala 40:28]
  assign PECross_12_multiply_io_input_io_actOut_ready = PECross_13_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_12_multiply_io_input_io_weiOut_ready = PECross_28_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_13_clock = clock;
  assign PECross_13_reset = rst;
  assign PECross_13_multiply_io_input_io_sumIn_valid = PECross_12_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_13_multiply_io_input_io_sumIn_bits_x_0 = PECross_12_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_13_multiply_io_input_io_sumIn_bits_last = PECross_12_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_13_multiply_io_input_io_sumOut_ready = PECross_14_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_13_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_13_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_13_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_13_multiply_io_input_io_actIn_valid = PECross_12_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_13_multiply_io_input_io_actIn_bits_x_0 = PECross_12_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_13_multiply_io_input_io_actIn_bits_last = PECross_12_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_13_multiply_io_input_io_weiIn_valid = io_weiIn_13_valid; // @[mac.scala 40:28]
  assign PECross_13_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_13_bits_x_0; // @[mac.scala 40:28]
  assign PECross_13_multiply_io_input_io_weiIn_bits_last = io_weiIn_13_bits_last; // @[mac.scala 40:28]
  assign PECross_13_multiply_io_input_io_actOut_ready = PECross_14_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_13_multiply_io_input_io_weiOut_ready = PECross_29_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_14_clock = clock;
  assign PECross_14_reset = rst;
  assign PECross_14_multiply_io_input_io_sumIn_valid = PECross_13_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_14_multiply_io_input_io_sumIn_bits_x_0 = PECross_13_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_14_multiply_io_input_io_sumIn_bits_last = PECross_13_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_14_multiply_io_input_io_sumOut_ready = PECross_15_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_14_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_14_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_14_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_14_multiply_io_input_io_actIn_valid = PECross_13_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_14_multiply_io_input_io_actIn_bits_x_0 = PECross_13_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_14_multiply_io_input_io_actIn_bits_last = PECross_13_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_14_multiply_io_input_io_weiIn_valid = io_weiIn_14_valid; // @[mac.scala 40:28]
  assign PECross_14_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_14_bits_x_0; // @[mac.scala 40:28]
  assign PECross_14_multiply_io_input_io_weiIn_bits_last = io_weiIn_14_bits_last; // @[mac.scala 40:28]
  assign PECross_14_multiply_io_input_io_actOut_ready = PECross_15_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_14_multiply_io_input_io_weiOut_ready = PECross_30_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_15_clock = clock;
  assign PECross_15_reset = rst;
  assign PECross_15_multiply_io_input_io_sumIn_valid = PECross_14_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_15_multiply_io_input_io_sumIn_bits_x_0 = PECross_14_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_15_multiply_io_input_io_sumIn_bits_last = PECross_14_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_15_multiply_io_input_io_sumOut_ready = io_sumOut_0_ready; // @[mac.scala 45:29]
  assign PECross_15_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_15_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_15_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_15_multiply_io_input_io_actIn_valid = PECross_14_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_15_multiply_io_input_io_actIn_bits_x_0 = PECross_14_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_15_multiply_io_input_io_actIn_bits_last = PECross_14_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_15_multiply_io_input_io_weiIn_valid = io_weiIn_15_valid; // @[mac.scala 40:28]
  assign PECross_15_multiply_io_input_io_weiIn_bits_x_0 = io_weiIn_15_bits_x_0; // @[mac.scala 40:28]
  assign PECross_15_multiply_io_input_io_weiIn_bits_last = io_weiIn_15_bits_last; // @[mac.scala 40:28]
  assign PECross_15_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_15_multiply_io_input_io_weiOut_ready = PECross_31_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_16_clock = clock;
  assign PECross_16_reset = rst;
  assign PECross_16_multiply_io_input_io_sumIn_valid = io_sumIn_1_valid; // @[mac.scala 33:28]
  assign PECross_16_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_1_bits_x_0; // @[mac.scala 33:28]
  assign PECross_16_multiply_io_input_io_sumIn_bits_last = io_sumIn_1_bits_last; // @[mac.scala 33:28]
  assign PECross_16_multiply_io_input_io_sumOut_ready = PECross_17_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_16_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_16_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_16_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_16_multiply_io_input_io_actIn_valid = io_actIn_1_valid; // @[mac.scala 32:28]
  assign PECross_16_multiply_io_input_io_actIn_bits_x_0 = io_actIn_1_bits_x_0; // @[mac.scala 32:28]
  assign PECross_16_multiply_io_input_io_actIn_bits_last = io_actIn_1_bits_last; // @[mac.scala 32:28]
  assign PECross_16_multiply_io_input_io_weiIn_valid = PECross_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_16_multiply_io_input_io_weiIn_bits_x_0 = PECross_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_16_multiply_io_input_io_weiIn_bits_last = PECross_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_16_multiply_io_input_io_actOut_ready = PECross_17_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_16_multiply_io_input_io_weiOut_ready = PECross_32_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_17_clock = clock;
  assign PECross_17_reset = rst;
  assign PECross_17_multiply_io_input_io_sumIn_valid = PECross_16_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_17_multiply_io_input_io_sumIn_bits_x_0 = PECross_16_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_17_multiply_io_input_io_sumIn_bits_last = PECross_16_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_17_multiply_io_input_io_sumOut_ready = PECross_18_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_17_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_17_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_17_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_17_multiply_io_input_io_actIn_valid = PECross_16_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_17_multiply_io_input_io_actIn_bits_x_0 = PECross_16_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_17_multiply_io_input_io_actIn_bits_last = PECross_16_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_17_multiply_io_input_io_weiIn_valid = PECross_1_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_17_multiply_io_input_io_weiIn_bits_x_0 = PECross_1_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_17_multiply_io_input_io_weiIn_bits_last = PECross_1_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_17_multiply_io_input_io_actOut_ready = PECross_18_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_17_multiply_io_input_io_weiOut_ready = PECross_33_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_18_clock = clock;
  assign PECross_18_reset = rst;
  assign PECross_18_multiply_io_input_io_sumIn_valid = PECross_17_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_18_multiply_io_input_io_sumIn_bits_x_0 = PECross_17_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_18_multiply_io_input_io_sumIn_bits_last = PECross_17_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_18_multiply_io_input_io_sumOut_ready = PECross_19_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_18_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_18_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_18_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_18_multiply_io_input_io_actIn_valid = PECross_17_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_18_multiply_io_input_io_actIn_bits_x_0 = PECross_17_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_18_multiply_io_input_io_actIn_bits_last = PECross_17_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_18_multiply_io_input_io_weiIn_valid = PECross_2_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_18_multiply_io_input_io_weiIn_bits_x_0 = PECross_2_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_18_multiply_io_input_io_weiIn_bits_last = PECross_2_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_18_multiply_io_input_io_actOut_ready = PECross_19_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_18_multiply_io_input_io_weiOut_ready = PECross_34_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_19_clock = clock;
  assign PECross_19_reset = rst;
  assign PECross_19_multiply_io_input_io_sumIn_valid = PECross_18_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_19_multiply_io_input_io_sumIn_bits_x_0 = PECross_18_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_19_multiply_io_input_io_sumIn_bits_last = PECross_18_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_19_multiply_io_input_io_sumOut_ready = PECross_20_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_19_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_19_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_19_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_19_multiply_io_input_io_actIn_valid = PECross_18_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_19_multiply_io_input_io_actIn_bits_x_0 = PECross_18_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_19_multiply_io_input_io_actIn_bits_last = PECross_18_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_19_multiply_io_input_io_weiIn_valid = PECross_3_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_19_multiply_io_input_io_weiIn_bits_x_0 = PECross_3_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_19_multiply_io_input_io_weiIn_bits_last = PECross_3_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_19_multiply_io_input_io_actOut_ready = PECross_20_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_19_multiply_io_input_io_weiOut_ready = PECross_35_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_20_clock = clock;
  assign PECross_20_reset = rst;
  assign PECross_20_multiply_io_input_io_sumIn_valid = PECross_19_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_20_multiply_io_input_io_sumIn_bits_x_0 = PECross_19_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_20_multiply_io_input_io_sumIn_bits_last = PECross_19_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_20_multiply_io_input_io_sumOut_ready = PECross_21_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_20_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_20_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_20_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_20_multiply_io_input_io_actIn_valid = PECross_19_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_20_multiply_io_input_io_actIn_bits_x_0 = PECross_19_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_20_multiply_io_input_io_actIn_bits_last = PECross_19_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_20_multiply_io_input_io_weiIn_valid = PECross_4_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_20_multiply_io_input_io_weiIn_bits_x_0 = PECross_4_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_20_multiply_io_input_io_weiIn_bits_last = PECross_4_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_20_multiply_io_input_io_actOut_ready = PECross_21_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_20_multiply_io_input_io_weiOut_ready = PECross_36_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_21_clock = clock;
  assign PECross_21_reset = rst;
  assign PECross_21_multiply_io_input_io_sumIn_valid = PECross_20_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_21_multiply_io_input_io_sumIn_bits_x_0 = PECross_20_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_21_multiply_io_input_io_sumIn_bits_last = PECross_20_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_21_multiply_io_input_io_sumOut_ready = PECross_22_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_21_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_21_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_21_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_21_multiply_io_input_io_actIn_valid = PECross_20_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_21_multiply_io_input_io_actIn_bits_x_0 = PECross_20_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_21_multiply_io_input_io_actIn_bits_last = PECross_20_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_21_multiply_io_input_io_weiIn_valid = PECross_5_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_21_multiply_io_input_io_weiIn_bits_x_0 = PECross_5_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_21_multiply_io_input_io_weiIn_bits_last = PECross_5_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_21_multiply_io_input_io_actOut_ready = PECross_22_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_21_multiply_io_input_io_weiOut_ready = PECross_37_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_22_clock = clock;
  assign PECross_22_reset = rst;
  assign PECross_22_multiply_io_input_io_sumIn_valid = PECross_21_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_22_multiply_io_input_io_sumIn_bits_x_0 = PECross_21_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_22_multiply_io_input_io_sumIn_bits_last = PECross_21_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_22_multiply_io_input_io_sumOut_ready = PECross_23_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_22_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_22_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_22_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_22_multiply_io_input_io_actIn_valid = PECross_21_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_22_multiply_io_input_io_actIn_bits_x_0 = PECross_21_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_22_multiply_io_input_io_actIn_bits_last = PECross_21_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_22_multiply_io_input_io_weiIn_valid = PECross_6_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_22_multiply_io_input_io_weiIn_bits_x_0 = PECross_6_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_22_multiply_io_input_io_weiIn_bits_last = PECross_6_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_22_multiply_io_input_io_actOut_ready = PECross_23_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_22_multiply_io_input_io_weiOut_ready = PECross_38_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_23_clock = clock;
  assign PECross_23_reset = rst;
  assign PECross_23_multiply_io_input_io_sumIn_valid = PECross_22_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_23_multiply_io_input_io_sumIn_bits_x_0 = PECross_22_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_23_multiply_io_input_io_sumIn_bits_last = PECross_22_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_23_multiply_io_input_io_sumOut_ready = PECross_24_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_23_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_23_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_23_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_23_multiply_io_input_io_actIn_valid = PECross_22_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_23_multiply_io_input_io_actIn_bits_x_0 = PECross_22_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_23_multiply_io_input_io_actIn_bits_last = PECross_22_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_23_multiply_io_input_io_weiIn_valid = PECross_7_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_23_multiply_io_input_io_weiIn_bits_x_0 = PECross_7_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_23_multiply_io_input_io_weiIn_bits_last = PECross_7_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_23_multiply_io_input_io_actOut_ready = PECross_24_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_23_multiply_io_input_io_weiOut_ready = PECross_39_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_24_clock = clock;
  assign PECross_24_reset = rst;
  assign PECross_24_multiply_io_input_io_sumIn_valid = PECross_23_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_24_multiply_io_input_io_sumIn_bits_x_0 = PECross_23_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_24_multiply_io_input_io_sumIn_bits_last = PECross_23_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_24_multiply_io_input_io_sumOut_ready = PECross_25_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_24_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_24_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_24_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_24_multiply_io_input_io_actIn_valid = PECross_23_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_24_multiply_io_input_io_actIn_bits_x_0 = PECross_23_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_24_multiply_io_input_io_actIn_bits_last = PECross_23_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_24_multiply_io_input_io_weiIn_valid = PECross_8_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_24_multiply_io_input_io_weiIn_bits_x_0 = PECross_8_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_24_multiply_io_input_io_weiIn_bits_last = PECross_8_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_24_multiply_io_input_io_actOut_ready = PECross_25_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_24_multiply_io_input_io_weiOut_ready = PECross_40_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_25_clock = clock;
  assign PECross_25_reset = rst;
  assign PECross_25_multiply_io_input_io_sumIn_valid = PECross_24_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_25_multiply_io_input_io_sumIn_bits_x_0 = PECross_24_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_25_multiply_io_input_io_sumIn_bits_last = PECross_24_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_25_multiply_io_input_io_sumOut_ready = PECross_26_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_25_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_25_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_25_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_25_multiply_io_input_io_actIn_valid = PECross_24_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_25_multiply_io_input_io_actIn_bits_x_0 = PECross_24_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_25_multiply_io_input_io_actIn_bits_last = PECross_24_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_25_multiply_io_input_io_weiIn_valid = PECross_9_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_25_multiply_io_input_io_weiIn_bits_x_0 = PECross_9_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_25_multiply_io_input_io_weiIn_bits_last = PECross_9_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_25_multiply_io_input_io_actOut_ready = PECross_26_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_25_multiply_io_input_io_weiOut_ready = PECross_41_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_26_clock = clock;
  assign PECross_26_reset = rst;
  assign PECross_26_multiply_io_input_io_sumIn_valid = PECross_25_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_26_multiply_io_input_io_sumIn_bits_x_0 = PECross_25_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_26_multiply_io_input_io_sumIn_bits_last = PECross_25_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_26_multiply_io_input_io_sumOut_ready = PECross_27_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_26_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_26_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_26_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_26_multiply_io_input_io_actIn_valid = PECross_25_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_26_multiply_io_input_io_actIn_bits_x_0 = PECross_25_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_26_multiply_io_input_io_actIn_bits_last = PECross_25_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_26_multiply_io_input_io_weiIn_valid = PECross_10_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_26_multiply_io_input_io_weiIn_bits_x_0 = PECross_10_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_26_multiply_io_input_io_weiIn_bits_last = PECross_10_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_26_multiply_io_input_io_actOut_ready = PECross_27_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_26_multiply_io_input_io_weiOut_ready = PECross_42_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_27_clock = clock;
  assign PECross_27_reset = rst;
  assign PECross_27_multiply_io_input_io_sumIn_valid = PECross_26_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_27_multiply_io_input_io_sumIn_bits_x_0 = PECross_26_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_27_multiply_io_input_io_sumIn_bits_last = PECross_26_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_27_multiply_io_input_io_sumOut_ready = PECross_28_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_27_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_27_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_27_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_27_multiply_io_input_io_actIn_valid = PECross_26_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_27_multiply_io_input_io_actIn_bits_x_0 = PECross_26_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_27_multiply_io_input_io_actIn_bits_last = PECross_26_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_27_multiply_io_input_io_weiIn_valid = PECross_11_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_27_multiply_io_input_io_weiIn_bits_x_0 = PECross_11_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_27_multiply_io_input_io_weiIn_bits_last = PECross_11_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_27_multiply_io_input_io_actOut_ready = PECross_28_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_27_multiply_io_input_io_weiOut_ready = PECross_43_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_28_clock = clock;
  assign PECross_28_reset = rst;
  assign PECross_28_multiply_io_input_io_sumIn_valid = PECross_27_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_28_multiply_io_input_io_sumIn_bits_x_0 = PECross_27_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_28_multiply_io_input_io_sumIn_bits_last = PECross_27_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_28_multiply_io_input_io_sumOut_ready = PECross_29_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_28_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_28_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_28_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_28_multiply_io_input_io_actIn_valid = PECross_27_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_28_multiply_io_input_io_actIn_bits_x_0 = PECross_27_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_28_multiply_io_input_io_actIn_bits_last = PECross_27_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_28_multiply_io_input_io_weiIn_valid = PECross_12_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_28_multiply_io_input_io_weiIn_bits_x_0 = PECross_12_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_28_multiply_io_input_io_weiIn_bits_last = PECross_12_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_28_multiply_io_input_io_actOut_ready = PECross_29_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_28_multiply_io_input_io_weiOut_ready = PECross_44_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_29_clock = clock;
  assign PECross_29_reset = rst;
  assign PECross_29_multiply_io_input_io_sumIn_valid = PECross_28_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_29_multiply_io_input_io_sumIn_bits_x_0 = PECross_28_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_29_multiply_io_input_io_sumIn_bits_last = PECross_28_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_29_multiply_io_input_io_sumOut_ready = PECross_30_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_29_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_29_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_29_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_29_multiply_io_input_io_actIn_valid = PECross_28_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_29_multiply_io_input_io_actIn_bits_x_0 = PECross_28_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_29_multiply_io_input_io_actIn_bits_last = PECross_28_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_29_multiply_io_input_io_weiIn_valid = PECross_13_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_29_multiply_io_input_io_weiIn_bits_x_0 = PECross_13_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_29_multiply_io_input_io_weiIn_bits_last = PECross_13_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_29_multiply_io_input_io_actOut_ready = PECross_30_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_29_multiply_io_input_io_weiOut_ready = PECross_45_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_30_clock = clock;
  assign PECross_30_reset = rst;
  assign PECross_30_multiply_io_input_io_sumIn_valid = PECross_29_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_30_multiply_io_input_io_sumIn_bits_x_0 = PECross_29_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_30_multiply_io_input_io_sumIn_bits_last = PECross_29_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_30_multiply_io_input_io_sumOut_ready = PECross_31_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_30_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_30_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_30_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_30_multiply_io_input_io_actIn_valid = PECross_29_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_30_multiply_io_input_io_actIn_bits_x_0 = PECross_29_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_30_multiply_io_input_io_actIn_bits_last = PECross_29_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_30_multiply_io_input_io_weiIn_valid = PECross_14_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_30_multiply_io_input_io_weiIn_bits_x_0 = PECross_14_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_30_multiply_io_input_io_weiIn_bits_last = PECross_14_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_30_multiply_io_input_io_actOut_ready = PECross_31_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_30_multiply_io_input_io_weiOut_ready = PECross_46_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_31_clock = clock;
  assign PECross_31_reset = rst;
  assign PECross_31_multiply_io_input_io_sumIn_valid = PECross_30_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_31_multiply_io_input_io_sumIn_bits_x_0 = PECross_30_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_31_multiply_io_input_io_sumIn_bits_last = PECross_30_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_31_multiply_io_input_io_sumOut_ready = io_sumOut_1_ready; // @[mac.scala 45:29]
  assign PECross_31_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_31_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_31_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_31_multiply_io_input_io_actIn_valid = PECross_30_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_31_multiply_io_input_io_actIn_bits_x_0 = PECross_30_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_31_multiply_io_input_io_actIn_bits_last = PECross_30_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_31_multiply_io_input_io_weiIn_valid = PECross_15_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_31_multiply_io_input_io_weiIn_bits_x_0 = PECross_15_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_31_multiply_io_input_io_weiIn_bits_last = PECross_15_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_31_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_31_multiply_io_input_io_weiOut_ready = PECross_47_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_32_clock = clock;
  assign PECross_32_reset = rst;
  assign PECross_32_multiply_io_input_io_sumIn_valid = io_sumIn_2_valid; // @[mac.scala 33:28]
  assign PECross_32_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_2_bits_x_0; // @[mac.scala 33:28]
  assign PECross_32_multiply_io_input_io_sumIn_bits_last = io_sumIn_2_bits_last; // @[mac.scala 33:28]
  assign PECross_32_multiply_io_input_io_sumOut_ready = PECross_33_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_32_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_32_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_32_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_32_multiply_io_input_io_actIn_valid = io_actIn_2_valid; // @[mac.scala 32:28]
  assign PECross_32_multiply_io_input_io_actIn_bits_x_0 = io_actIn_2_bits_x_0; // @[mac.scala 32:28]
  assign PECross_32_multiply_io_input_io_actIn_bits_last = io_actIn_2_bits_last; // @[mac.scala 32:28]
  assign PECross_32_multiply_io_input_io_weiIn_valid = PECross_16_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_32_multiply_io_input_io_weiIn_bits_x_0 = PECross_16_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_32_multiply_io_input_io_weiIn_bits_last = PECross_16_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_32_multiply_io_input_io_actOut_ready = PECross_33_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_32_multiply_io_input_io_weiOut_ready = PECross_48_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_33_clock = clock;
  assign PECross_33_reset = rst;
  assign PECross_33_multiply_io_input_io_sumIn_valid = PECross_32_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_33_multiply_io_input_io_sumIn_bits_x_0 = PECross_32_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_33_multiply_io_input_io_sumIn_bits_last = PECross_32_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_33_multiply_io_input_io_sumOut_ready = PECross_34_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_33_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_33_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_33_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_33_multiply_io_input_io_actIn_valid = PECross_32_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_33_multiply_io_input_io_actIn_bits_x_0 = PECross_32_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_33_multiply_io_input_io_actIn_bits_last = PECross_32_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_33_multiply_io_input_io_weiIn_valid = PECross_17_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_33_multiply_io_input_io_weiIn_bits_x_0 = PECross_17_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_33_multiply_io_input_io_weiIn_bits_last = PECross_17_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_33_multiply_io_input_io_actOut_ready = PECross_34_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_33_multiply_io_input_io_weiOut_ready = PECross_49_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_34_clock = clock;
  assign PECross_34_reset = rst;
  assign PECross_34_multiply_io_input_io_sumIn_valid = PECross_33_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_34_multiply_io_input_io_sumIn_bits_x_0 = PECross_33_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_34_multiply_io_input_io_sumIn_bits_last = PECross_33_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_34_multiply_io_input_io_sumOut_ready = PECross_35_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_34_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_34_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_34_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_34_multiply_io_input_io_actIn_valid = PECross_33_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_34_multiply_io_input_io_actIn_bits_x_0 = PECross_33_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_34_multiply_io_input_io_actIn_bits_last = PECross_33_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_34_multiply_io_input_io_weiIn_valid = PECross_18_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_34_multiply_io_input_io_weiIn_bits_x_0 = PECross_18_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_34_multiply_io_input_io_weiIn_bits_last = PECross_18_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_34_multiply_io_input_io_actOut_ready = PECross_35_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_34_multiply_io_input_io_weiOut_ready = PECross_50_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_35_clock = clock;
  assign PECross_35_reset = rst;
  assign PECross_35_multiply_io_input_io_sumIn_valid = PECross_34_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_35_multiply_io_input_io_sumIn_bits_x_0 = PECross_34_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_35_multiply_io_input_io_sumIn_bits_last = PECross_34_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_35_multiply_io_input_io_sumOut_ready = PECross_36_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_35_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_35_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_35_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_35_multiply_io_input_io_actIn_valid = PECross_34_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_35_multiply_io_input_io_actIn_bits_x_0 = PECross_34_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_35_multiply_io_input_io_actIn_bits_last = PECross_34_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_35_multiply_io_input_io_weiIn_valid = PECross_19_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_35_multiply_io_input_io_weiIn_bits_x_0 = PECross_19_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_35_multiply_io_input_io_weiIn_bits_last = PECross_19_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_35_multiply_io_input_io_actOut_ready = PECross_36_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_35_multiply_io_input_io_weiOut_ready = PECross_51_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_36_clock = clock;
  assign PECross_36_reset = rst;
  assign PECross_36_multiply_io_input_io_sumIn_valid = PECross_35_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_36_multiply_io_input_io_sumIn_bits_x_0 = PECross_35_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_36_multiply_io_input_io_sumIn_bits_last = PECross_35_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_36_multiply_io_input_io_sumOut_ready = PECross_37_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_36_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_36_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_36_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_36_multiply_io_input_io_actIn_valid = PECross_35_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_36_multiply_io_input_io_actIn_bits_x_0 = PECross_35_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_36_multiply_io_input_io_actIn_bits_last = PECross_35_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_36_multiply_io_input_io_weiIn_valid = PECross_20_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_36_multiply_io_input_io_weiIn_bits_x_0 = PECross_20_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_36_multiply_io_input_io_weiIn_bits_last = PECross_20_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_36_multiply_io_input_io_actOut_ready = PECross_37_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_36_multiply_io_input_io_weiOut_ready = PECross_52_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_37_clock = clock;
  assign PECross_37_reset = rst;
  assign PECross_37_multiply_io_input_io_sumIn_valid = PECross_36_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_37_multiply_io_input_io_sumIn_bits_x_0 = PECross_36_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_37_multiply_io_input_io_sumIn_bits_last = PECross_36_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_37_multiply_io_input_io_sumOut_ready = PECross_38_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_37_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_37_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_37_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_37_multiply_io_input_io_actIn_valid = PECross_36_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_37_multiply_io_input_io_actIn_bits_x_0 = PECross_36_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_37_multiply_io_input_io_actIn_bits_last = PECross_36_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_37_multiply_io_input_io_weiIn_valid = PECross_21_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_37_multiply_io_input_io_weiIn_bits_x_0 = PECross_21_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_37_multiply_io_input_io_weiIn_bits_last = PECross_21_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_37_multiply_io_input_io_actOut_ready = PECross_38_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_37_multiply_io_input_io_weiOut_ready = PECross_53_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_38_clock = clock;
  assign PECross_38_reset = rst;
  assign PECross_38_multiply_io_input_io_sumIn_valid = PECross_37_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_38_multiply_io_input_io_sumIn_bits_x_0 = PECross_37_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_38_multiply_io_input_io_sumIn_bits_last = PECross_37_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_38_multiply_io_input_io_sumOut_ready = PECross_39_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_38_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_38_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_38_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_38_multiply_io_input_io_actIn_valid = PECross_37_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_38_multiply_io_input_io_actIn_bits_x_0 = PECross_37_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_38_multiply_io_input_io_actIn_bits_last = PECross_37_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_38_multiply_io_input_io_weiIn_valid = PECross_22_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_38_multiply_io_input_io_weiIn_bits_x_0 = PECross_22_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_38_multiply_io_input_io_weiIn_bits_last = PECross_22_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_38_multiply_io_input_io_actOut_ready = PECross_39_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_38_multiply_io_input_io_weiOut_ready = PECross_54_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_39_clock = clock;
  assign PECross_39_reset = rst;
  assign PECross_39_multiply_io_input_io_sumIn_valid = PECross_38_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_39_multiply_io_input_io_sumIn_bits_x_0 = PECross_38_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_39_multiply_io_input_io_sumIn_bits_last = PECross_38_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_39_multiply_io_input_io_sumOut_ready = PECross_40_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_39_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_39_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_39_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_39_multiply_io_input_io_actIn_valid = PECross_38_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_39_multiply_io_input_io_actIn_bits_x_0 = PECross_38_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_39_multiply_io_input_io_actIn_bits_last = PECross_38_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_39_multiply_io_input_io_weiIn_valid = PECross_23_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_39_multiply_io_input_io_weiIn_bits_x_0 = PECross_23_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_39_multiply_io_input_io_weiIn_bits_last = PECross_23_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_39_multiply_io_input_io_actOut_ready = PECross_40_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_39_multiply_io_input_io_weiOut_ready = PECross_55_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_40_clock = clock;
  assign PECross_40_reset = rst;
  assign PECross_40_multiply_io_input_io_sumIn_valid = PECross_39_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_40_multiply_io_input_io_sumIn_bits_x_0 = PECross_39_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_40_multiply_io_input_io_sumIn_bits_last = PECross_39_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_40_multiply_io_input_io_sumOut_ready = PECross_41_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_40_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_40_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_40_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_40_multiply_io_input_io_actIn_valid = PECross_39_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_40_multiply_io_input_io_actIn_bits_x_0 = PECross_39_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_40_multiply_io_input_io_actIn_bits_last = PECross_39_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_40_multiply_io_input_io_weiIn_valid = PECross_24_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_40_multiply_io_input_io_weiIn_bits_x_0 = PECross_24_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_40_multiply_io_input_io_weiIn_bits_last = PECross_24_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_40_multiply_io_input_io_actOut_ready = PECross_41_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_40_multiply_io_input_io_weiOut_ready = PECross_56_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_41_clock = clock;
  assign PECross_41_reset = rst;
  assign PECross_41_multiply_io_input_io_sumIn_valid = PECross_40_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_41_multiply_io_input_io_sumIn_bits_x_0 = PECross_40_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_41_multiply_io_input_io_sumIn_bits_last = PECross_40_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_41_multiply_io_input_io_sumOut_ready = PECross_42_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_41_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_41_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_41_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_41_multiply_io_input_io_actIn_valid = PECross_40_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_41_multiply_io_input_io_actIn_bits_x_0 = PECross_40_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_41_multiply_io_input_io_actIn_bits_last = PECross_40_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_41_multiply_io_input_io_weiIn_valid = PECross_25_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_41_multiply_io_input_io_weiIn_bits_x_0 = PECross_25_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_41_multiply_io_input_io_weiIn_bits_last = PECross_25_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_41_multiply_io_input_io_actOut_ready = PECross_42_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_41_multiply_io_input_io_weiOut_ready = PECross_57_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_42_clock = clock;
  assign PECross_42_reset = rst;
  assign PECross_42_multiply_io_input_io_sumIn_valid = PECross_41_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_42_multiply_io_input_io_sumIn_bits_x_0 = PECross_41_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_42_multiply_io_input_io_sumIn_bits_last = PECross_41_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_42_multiply_io_input_io_sumOut_ready = PECross_43_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_42_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_42_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_42_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_42_multiply_io_input_io_actIn_valid = PECross_41_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_42_multiply_io_input_io_actIn_bits_x_0 = PECross_41_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_42_multiply_io_input_io_actIn_bits_last = PECross_41_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_42_multiply_io_input_io_weiIn_valid = PECross_26_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_42_multiply_io_input_io_weiIn_bits_x_0 = PECross_26_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_42_multiply_io_input_io_weiIn_bits_last = PECross_26_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_42_multiply_io_input_io_actOut_ready = PECross_43_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_42_multiply_io_input_io_weiOut_ready = PECross_58_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_43_clock = clock;
  assign PECross_43_reset = rst;
  assign PECross_43_multiply_io_input_io_sumIn_valid = PECross_42_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_43_multiply_io_input_io_sumIn_bits_x_0 = PECross_42_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_43_multiply_io_input_io_sumIn_bits_last = PECross_42_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_43_multiply_io_input_io_sumOut_ready = PECross_44_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_43_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_43_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_43_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_43_multiply_io_input_io_actIn_valid = PECross_42_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_43_multiply_io_input_io_actIn_bits_x_0 = PECross_42_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_43_multiply_io_input_io_actIn_bits_last = PECross_42_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_43_multiply_io_input_io_weiIn_valid = PECross_27_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_43_multiply_io_input_io_weiIn_bits_x_0 = PECross_27_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_43_multiply_io_input_io_weiIn_bits_last = PECross_27_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_43_multiply_io_input_io_actOut_ready = PECross_44_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_43_multiply_io_input_io_weiOut_ready = PECross_59_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_44_clock = clock;
  assign PECross_44_reset = rst;
  assign PECross_44_multiply_io_input_io_sumIn_valid = PECross_43_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_44_multiply_io_input_io_sumIn_bits_x_0 = PECross_43_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_44_multiply_io_input_io_sumIn_bits_last = PECross_43_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_44_multiply_io_input_io_sumOut_ready = PECross_45_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_44_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_44_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_44_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_44_multiply_io_input_io_actIn_valid = PECross_43_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_44_multiply_io_input_io_actIn_bits_x_0 = PECross_43_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_44_multiply_io_input_io_actIn_bits_last = PECross_43_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_44_multiply_io_input_io_weiIn_valid = PECross_28_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_44_multiply_io_input_io_weiIn_bits_x_0 = PECross_28_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_44_multiply_io_input_io_weiIn_bits_last = PECross_28_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_44_multiply_io_input_io_actOut_ready = PECross_45_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_44_multiply_io_input_io_weiOut_ready = PECross_60_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_45_clock = clock;
  assign PECross_45_reset = rst;
  assign PECross_45_multiply_io_input_io_sumIn_valid = PECross_44_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_45_multiply_io_input_io_sumIn_bits_x_0 = PECross_44_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_45_multiply_io_input_io_sumIn_bits_last = PECross_44_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_45_multiply_io_input_io_sumOut_ready = PECross_46_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_45_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_45_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_45_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_45_multiply_io_input_io_actIn_valid = PECross_44_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_45_multiply_io_input_io_actIn_bits_x_0 = PECross_44_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_45_multiply_io_input_io_actIn_bits_last = PECross_44_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_45_multiply_io_input_io_weiIn_valid = PECross_29_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_45_multiply_io_input_io_weiIn_bits_x_0 = PECross_29_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_45_multiply_io_input_io_weiIn_bits_last = PECross_29_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_45_multiply_io_input_io_actOut_ready = PECross_46_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_45_multiply_io_input_io_weiOut_ready = PECross_61_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_46_clock = clock;
  assign PECross_46_reset = rst;
  assign PECross_46_multiply_io_input_io_sumIn_valid = PECross_45_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_46_multiply_io_input_io_sumIn_bits_x_0 = PECross_45_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_46_multiply_io_input_io_sumIn_bits_last = PECross_45_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_46_multiply_io_input_io_sumOut_ready = PECross_47_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_46_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_46_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_46_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_46_multiply_io_input_io_actIn_valid = PECross_45_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_46_multiply_io_input_io_actIn_bits_x_0 = PECross_45_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_46_multiply_io_input_io_actIn_bits_last = PECross_45_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_46_multiply_io_input_io_weiIn_valid = PECross_30_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_46_multiply_io_input_io_weiIn_bits_x_0 = PECross_30_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_46_multiply_io_input_io_weiIn_bits_last = PECross_30_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_46_multiply_io_input_io_actOut_ready = PECross_47_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_46_multiply_io_input_io_weiOut_ready = PECross_62_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_47_clock = clock;
  assign PECross_47_reset = rst;
  assign PECross_47_multiply_io_input_io_sumIn_valid = PECross_46_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_47_multiply_io_input_io_sumIn_bits_x_0 = PECross_46_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_47_multiply_io_input_io_sumIn_bits_last = PECross_46_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_47_multiply_io_input_io_sumOut_ready = io_sumOut_2_ready; // @[mac.scala 45:29]
  assign PECross_47_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_47_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_47_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_47_multiply_io_input_io_actIn_valid = PECross_46_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_47_multiply_io_input_io_actIn_bits_x_0 = PECross_46_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_47_multiply_io_input_io_actIn_bits_last = PECross_46_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_47_multiply_io_input_io_weiIn_valid = PECross_31_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_47_multiply_io_input_io_weiIn_bits_x_0 = PECross_31_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_47_multiply_io_input_io_weiIn_bits_last = PECross_31_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_47_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_47_multiply_io_input_io_weiOut_ready = PECross_63_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_48_clock = clock;
  assign PECross_48_reset = rst;
  assign PECross_48_multiply_io_input_io_sumIn_valid = io_sumIn_3_valid; // @[mac.scala 33:28]
  assign PECross_48_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_3_bits_x_0; // @[mac.scala 33:28]
  assign PECross_48_multiply_io_input_io_sumIn_bits_last = io_sumIn_3_bits_last; // @[mac.scala 33:28]
  assign PECross_48_multiply_io_input_io_sumOut_ready = PECross_49_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_48_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_48_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_48_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_48_multiply_io_input_io_actIn_valid = io_actIn_3_valid; // @[mac.scala 32:28]
  assign PECross_48_multiply_io_input_io_actIn_bits_x_0 = io_actIn_3_bits_x_0; // @[mac.scala 32:28]
  assign PECross_48_multiply_io_input_io_actIn_bits_last = io_actIn_3_bits_last; // @[mac.scala 32:28]
  assign PECross_48_multiply_io_input_io_weiIn_valid = PECross_32_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_48_multiply_io_input_io_weiIn_bits_x_0 = PECross_32_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_48_multiply_io_input_io_weiIn_bits_last = PECross_32_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_48_multiply_io_input_io_actOut_ready = PECross_49_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_48_multiply_io_input_io_weiOut_ready = PECross_64_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_49_clock = clock;
  assign PECross_49_reset = rst;
  assign PECross_49_multiply_io_input_io_sumIn_valid = PECross_48_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_49_multiply_io_input_io_sumIn_bits_x_0 = PECross_48_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_49_multiply_io_input_io_sumIn_bits_last = PECross_48_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_49_multiply_io_input_io_sumOut_ready = PECross_50_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_49_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_49_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_49_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_49_multiply_io_input_io_actIn_valid = PECross_48_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_49_multiply_io_input_io_actIn_bits_x_0 = PECross_48_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_49_multiply_io_input_io_actIn_bits_last = PECross_48_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_49_multiply_io_input_io_weiIn_valid = PECross_33_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_49_multiply_io_input_io_weiIn_bits_x_0 = PECross_33_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_49_multiply_io_input_io_weiIn_bits_last = PECross_33_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_49_multiply_io_input_io_actOut_ready = PECross_50_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_49_multiply_io_input_io_weiOut_ready = PECross_65_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_50_clock = clock;
  assign PECross_50_reset = rst;
  assign PECross_50_multiply_io_input_io_sumIn_valid = PECross_49_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_50_multiply_io_input_io_sumIn_bits_x_0 = PECross_49_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_50_multiply_io_input_io_sumIn_bits_last = PECross_49_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_50_multiply_io_input_io_sumOut_ready = PECross_51_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_50_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_50_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_50_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_50_multiply_io_input_io_actIn_valid = PECross_49_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_50_multiply_io_input_io_actIn_bits_x_0 = PECross_49_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_50_multiply_io_input_io_actIn_bits_last = PECross_49_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_50_multiply_io_input_io_weiIn_valid = PECross_34_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_50_multiply_io_input_io_weiIn_bits_x_0 = PECross_34_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_50_multiply_io_input_io_weiIn_bits_last = PECross_34_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_50_multiply_io_input_io_actOut_ready = PECross_51_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_50_multiply_io_input_io_weiOut_ready = PECross_66_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_51_clock = clock;
  assign PECross_51_reset = rst;
  assign PECross_51_multiply_io_input_io_sumIn_valid = PECross_50_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_51_multiply_io_input_io_sumIn_bits_x_0 = PECross_50_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_51_multiply_io_input_io_sumIn_bits_last = PECross_50_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_51_multiply_io_input_io_sumOut_ready = PECross_52_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_51_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_51_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_51_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_51_multiply_io_input_io_actIn_valid = PECross_50_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_51_multiply_io_input_io_actIn_bits_x_0 = PECross_50_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_51_multiply_io_input_io_actIn_bits_last = PECross_50_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_51_multiply_io_input_io_weiIn_valid = PECross_35_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_51_multiply_io_input_io_weiIn_bits_x_0 = PECross_35_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_51_multiply_io_input_io_weiIn_bits_last = PECross_35_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_51_multiply_io_input_io_actOut_ready = PECross_52_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_51_multiply_io_input_io_weiOut_ready = PECross_67_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_52_clock = clock;
  assign PECross_52_reset = rst;
  assign PECross_52_multiply_io_input_io_sumIn_valid = PECross_51_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_52_multiply_io_input_io_sumIn_bits_x_0 = PECross_51_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_52_multiply_io_input_io_sumIn_bits_last = PECross_51_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_52_multiply_io_input_io_sumOut_ready = PECross_53_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_52_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_52_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_52_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_52_multiply_io_input_io_actIn_valid = PECross_51_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_52_multiply_io_input_io_actIn_bits_x_0 = PECross_51_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_52_multiply_io_input_io_actIn_bits_last = PECross_51_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_52_multiply_io_input_io_weiIn_valid = PECross_36_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_52_multiply_io_input_io_weiIn_bits_x_0 = PECross_36_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_52_multiply_io_input_io_weiIn_bits_last = PECross_36_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_52_multiply_io_input_io_actOut_ready = PECross_53_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_52_multiply_io_input_io_weiOut_ready = PECross_68_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_53_clock = clock;
  assign PECross_53_reset = rst;
  assign PECross_53_multiply_io_input_io_sumIn_valid = PECross_52_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_53_multiply_io_input_io_sumIn_bits_x_0 = PECross_52_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_53_multiply_io_input_io_sumIn_bits_last = PECross_52_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_53_multiply_io_input_io_sumOut_ready = PECross_54_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_53_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_53_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_53_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_53_multiply_io_input_io_actIn_valid = PECross_52_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_53_multiply_io_input_io_actIn_bits_x_0 = PECross_52_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_53_multiply_io_input_io_actIn_bits_last = PECross_52_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_53_multiply_io_input_io_weiIn_valid = PECross_37_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_53_multiply_io_input_io_weiIn_bits_x_0 = PECross_37_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_53_multiply_io_input_io_weiIn_bits_last = PECross_37_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_53_multiply_io_input_io_actOut_ready = PECross_54_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_53_multiply_io_input_io_weiOut_ready = PECross_69_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_54_clock = clock;
  assign PECross_54_reset = rst;
  assign PECross_54_multiply_io_input_io_sumIn_valid = PECross_53_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_54_multiply_io_input_io_sumIn_bits_x_0 = PECross_53_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_54_multiply_io_input_io_sumIn_bits_last = PECross_53_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_54_multiply_io_input_io_sumOut_ready = PECross_55_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_54_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_54_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_54_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_54_multiply_io_input_io_actIn_valid = PECross_53_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_54_multiply_io_input_io_actIn_bits_x_0 = PECross_53_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_54_multiply_io_input_io_actIn_bits_last = PECross_53_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_54_multiply_io_input_io_weiIn_valid = PECross_38_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_54_multiply_io_input_io_weiIn_bits_x_0 = PECross_38_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_54_multiply_io_input_io_weiIn_bits_last = PECross_38_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_54_multiply_io_input_io_actOut_ready = PECross_55_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_54_multiply_io_input_io_weiOut_ready = PECross_70_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_55_clock = clock;
  assign PECross_55_reset = rst;
  assign PECross_55_multiply_io_input_io_sumIn_valid = PECross_54_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_55_multiply_io_input_io_sumIn_bits_x_0 = PECross_54_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_55_multiply_io_input_io_sumIn_bits_last = PECross_54_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_55_multiply_io_input_io_sumOut_ready = PECross_56_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_55_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_55_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_55_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_55_multiply_io_input_io_actIn_valid = PECross_54_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_55_multiply_io_input_io_actIn_bits_x_0 = PECross_54_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_55_multiply_io_input_io_actIn_bits_last = PECross_54_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_55_multiply_io_input_io_weiIn_valid = PECross_39_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_55_multiply_io_input_io_weiIn_bits_x_0 = PECross_39_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_55_multiply_io_input_io_weiIn_bits_last = PECross_39_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_55_multiply_io_input_io_actOut_ready = PECross_56_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_55_multiply_io_input_io_weiOut_ready = PECross_71_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_56_clock = clock;
  assign PECross_56_reset = rst;
  assign PECross_56_multiply_io_input_io_sumIn_valid = PECross_55_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_56_multiply_io_input_io_sumIn_bits_x_0 = PECross_55_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_56_multiply_io_input_io_sumIn_bits_last = PECross_55_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_56_multiply_io_input_io_sumOut_ready = PECross_57_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_56_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_56_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_56_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_56_multiply_io_input_io_actIn_valid = PECross_55_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_56_multiply_io_input_io_actIn_bits_x_0 = PECross_55_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_56_multiply_io_input_io_actIn_bits_last = PECross_55_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_56_multiply_io_input_io_weiIn_valid = PECross_40_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_56_multiply_io_input_io_weiIn_bits_x_0 = PECross_40_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_56_multiply_io_input_io_weiIn_bits_last = PECross_40_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_56_multiply_io_input_io_actOut_ready = PECross_57_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_56_multiply_io_input_io_weiOut_ready = PECross_72_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_57_clock = clock;
  assign PECross_57_reset = rst;
  assign PECross_57_multiply_io_input_io_sumIn_valid = PECross_56_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_57_multiply_io_input_io_sumIn_bits_x_0 = PECross_56_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_57_multiply_io_input_io_sumIn_bits_last = PECross_56_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_57_multiply_io_input_io_sumOut_ready = PECross_58_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_57_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_57_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_57_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_57_multiply_io_input_io_actIn_valid = PECross_56_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_57_multiply_io_input_io_actIn_bits_x_0 = PECross_56_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_57_multiply_io_input_io_actIn_bits_last = PECross_56_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_57_multiply_io_input_io_weiIn_valid = PECross_41_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_57_multiply_io_input_io_weiIn_bits_x_0 = PECross_41_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_57_multiply_io_input_io_weiIn_bits_last = PECross_41_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_57_multiply_io_input_io_actOut_ready = PECross_58_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_57_multiply_io_input_io_weiOut_ready = PECross_73_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_58_clock = clock;
  assign PECross_58_reset = rst;
  assign PECross_58_multiply_io_input_io_sumIn_valid = PECross_57_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_58_multiply_io_input_io_sumIn_bits_x_0 = PECross_57_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_58_multiply_io_input_io_sumIn_bits_last = PECross_57_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_58_multiply_io_input_io_sumOut_ready = PECross_59_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_58_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_58_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_58_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_58_multiply_io_input_io_actIn_valid = PECross_57_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_58_multiply_io_input_io_actIn_bits_x_0 = PECross_57_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_58_multiply_io_input_io_actIn_bits_last = PECross_57_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_58_multiply_io_input_io_weiIn_valid = PECross_42_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_58_multiply_io_input_io_weiIn_bits_x_0 = PECross_42_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_58_multiply_io_input_io_weiIn_bits_last = PECross_42_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_58_multiply_io_input_io_actOut_ready = PECross_59_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_58_multiply_io_input_io_weiOut_ready = PECross_74_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_59_clock = clock;
  assign PECross_59_reset = rst;
  assign PECross_59_multiply_io_input_io_sumIn_valid = PECross_58_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_59_multiply_io_input_io_sumIn_bits_x_0 = PECross_58_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_59_multiply_io_input_io_sumIn_bits_last = PECross_58_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_59_multiply_io_input_io_sumOut_ready = PECross_60_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_59_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_59_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_59_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_59_multiply_io_input_io_actIn_valid = PECross_58_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_59_multiply_io_input_io_actIn_bits_x_0 = PECross_58_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_59_multiply_io_input_io_actIn_bits_last = PECross_58_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_59_multiply_io_input_io_weiIn_valid = PECross_43_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_59_multiply_io_input_io_weiIn_bits_x_0 = PECross_43_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_59_multiply_io_input_io_weiIn_bits_last = PECross_43_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_59_multiply_io_input_io_actOut_ready = PECross_60_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_59_multiply_io_input_io_weiOut_ready = PECross_75_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_60_clock = clock;
  assign PECross_60_reset = rst;
  assign PECross_60_multiply_io_input_io_sumIn_valid = PECross_59_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_60_multiply_io_input_io_sumIn_bits_x_0 = PECross_59_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_60_multiply_io_input_io_sumIn_bits_last = PECross_59_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_60_multiply_io_input_io_sumOut_ready = PECross_61_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_60_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_60_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_60_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_60_multiply_io_input_io_actIn_valid = PECross_59_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_60_multiply_io_input_io_actIn_bits_x_0 = PECross_59_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_60_multiply_io_input_io_actIn_bits_last = PECross_59_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_60_multiply_io_input_io_weiIn_valid = PECross_44_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_60_multiply_io_input_io_weiIn_bits_x_0 = PECross_44_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_60_multiply_io_input_io_weiIn_bits_last = PECross_44_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_60_multiply_io_input_io_actOut_ready = PECross_61_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_60_multiply_io_input_io_weiOut_ready = PECross_76_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_61_clock = clock;
  assign PECross_61_reset = rst;
  assign PECross_61_multiply_io_input_io_sumIn_valid = PECross_60_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_61_multiply_io_input_io_sumIn_bits_x_0 = PECross_60_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_61_multiply_io_input_io_sumIn_bits_last = PECross_60_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_61_multiply_io_input_io_sumOut_ready = PECross_62_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_61_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_61_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_61_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_61_multiply_io_input_io_actIn_valid = PECross_60_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_61_multiply_io_input_io_actIn_bits_x_0 = PECross_60_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_61_multiply_io_input_io_actIn_bits_last = PECross_60_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_61_multiply_io_input_io_weiIn_valid = PECross_45_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_61_multiply_io_input_io_weiIn_bits_x_0 = PECross_45_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_61_multiply_io_input_io_weiIn_bits_last = PECross_45_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_61_multiply_io_input_io_actOut_ready = PECross_62_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_61_multiply_io_input_io_weiOut_ready = PECross_77_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_62_clock = clock;
  assign PECross_62_reset = rst;
  assign PECross_62_multiply_io_input_io_sumIn_valid = PECross_61_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_62_multiply_io_input_io_sumIn_bits_x_0 = PECross_61_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_62_multiply_io_input_io_sumIn_bits_last = PECross_61_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_62_multiply_io_input_io_sumOut_ready = PECross_63_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_62_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_62_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_62_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_62_multiply_io_input_io_actIn_valid = PECross_61_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_62_multiply_io_input_io_actIn_bits_x_0 = PECross_61_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_62_multiply_io_input_io_actIn_bits_last = PECross_61_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_62_multiply_io_input_io_weiIn_valid = PECross_46_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_62_multiply_io_input_io_weiIn_bits_x_0 = PECross_46_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_62_multiply_io_input_io_weiIn_bits_last = PECross_46_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_62_multiply_io_input_io_actOut_ready = PECross_63_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_62_multiply_io_input_io_weiOut_ready = PECross_78_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_63_clock = clock;
  assign PECross_63_reset = rst;
  assign PECross_63_multiply_io_input_io_sumIn_valid = PECross_62_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_63_multiply_io_input_io_sumIn_bits_x_0 = PECross_62_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_63_multiply_io_input_io_sumIn_bits_last = PECross_62_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_63_multiply_io_input_io_sumOut_ready = io_sumOut_3_ready; // @[mac.scala 45:29]
  assign PECross_63_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_63_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_63_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_63_multiply_io_input_io_actIn_valid = PECross_62_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_63_multiply_io_input_io_actIn_bits_x_0 = PECross_62_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_63_multiply_io_input_io_actIn_bits_last = PECross_62_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_63_multiply_io_input_io_weiIn_valid = PECross_47_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_63_multiply_io_input_io_weiIn_bits_x_0 = PECross_47_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_63_multiply_io_input_io_weiIn_bits_last = PECross_47_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_63_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_63_multiply_io_input_io_weiOut_ready = PECross_79_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_64_clock = clock;
  assign PECross_64_reset = rst;
  assign PECross_64_multiply_io_input_io_sumIn_valid = io_sumIn_4_valid; // @[mac.scala 33:28]
  assign PECross_64_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_4_bits_x_0; // @[mac.scala 33:28]
  assign PECross_64_multiply_io_input_io_sumIn_bits_last = io_sumIn_4_bits_last; // @[mac.scala 33:28]
  assign PECross_64_multiply_io_input_io_sumOut_ready = PECross_65_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_64_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_64_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_64_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_64_multiply_io_input_io_actIn_valid = io_actIn_4_valid; // @[mac.scala 32:28]
  assign PECross_64_multiply_io_input_io_actIn_bits_x_0 = io_actIn_4_bits_x_0; // @[mac.scala 32:28]
  assign PECross_64_multiply_io_input_io_actIn_bits_last = io_actIn_4_bits_last; // @[mac.scala 32:28]
  assign PECross_64_multiply_io_input_io_weiIn_valid = PECross_48_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_64_multiply_io_input_io_weiIn_bits_x_0 = PECross_48_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_64_multiply_io_input_io_weiIn_bits_last = PECross_48_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_64_multiply_io_input_io_actOut_ready = PECross_65_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_64_multiply_io_input_io_weiOut_ready = PECross_80_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_65_clock = clock;
  assign PECross_65_reset = rst;
  assign PECross_65_multiply_io_input_io_sumIn_valid = PECross_64_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_65_multiply_io_input_io_sumIn_bits_x_0 = PECross_64_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_65_multiply_io_input_io_sumIn_bits_last = PECross_64_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_65_multiply_io_input_io_sumOut_ready = PECross_66_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_65_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_65_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_65_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_65_multiply_io_input_io_actIn_valid = PECross_64_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_65_multiply_io_input_io_actIn_bits_x_0 = PECross_64_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_65_multiply_io_input_io_actIn_bits_last = PECross_64_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_65_multiply_io_input_io_weiIn_valid = PECross_49_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_65_multiply_io_input_io_weiIn_bits_x_0 = PECross_49_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_65_multiply_io_input_io_weiIn_bits_last = PECross_49_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_65_multiply_io_input_io_actOut_ready = PECross_66_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_65_multiply_io_input_io_weiOut_ready = PECross_81_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_66_clock = clock;
  assign PECross_66_reset = rst;
  assign PECross_66_multiply_io_input_io_sumIn_valid = PECross_65_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_66_multiply_io_input_io_sumIn_bits_x_0 = PECross_65_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_66_multiply_io_input_io_sumIn_bits_last = PECross_65_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_66_multiply_io_input_io_sumOut_ready = PECross_67_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_66_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_66_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_66_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_66_multiply_io_input_io_actIn_valid = PECross_65_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_66_multiply_io_input_io_actIn_bits_x_0 = PECross_65_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_66_multiply_io_input_io_actIn_bits_last = PECross_65_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_66_multiply_io_input_io_weiIn_valid = PECross_50_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_66_multiply_io_input_io_weiIn_bits_x_0 = PECross_50_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_66_multiply_io_input_io_weiIn_bits_last = PECross_50_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_66_multiply_io_input_io_actOut_ready = PECross_67_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_66_multiply_io_input_io_weiOut_ready = PECross_82_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_67_clock = clock;
  assign PECross_67_reset = rst;
  assign PECross_67_multiply_io_input_io_sumIn_valid = PECross_66_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_67_multiply_io_input_io_sumIn_bits_x_0 = PECross_66_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_67_multiply_io_input_io_sumIn_bits_last = PECross_66_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_67_multiply_io_input_io_sumOut_ready = PECross_68_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_67_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_67_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_67_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_67_multiply_io_input_io_actIn_valid = PECross_66_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_67_multiply_io_input_io_actIn_bits_x_0 = PECross_66_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_67_multiply_io_input_io_actIn_bits_last = PECross_66_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_67_multiply_io_input_io_weiIn_valid = PECross_51_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_67_multiply_io_input_io_weiIn_bits_x_0 = PECross_51_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_67_multiply_io_input_io_weiIn_bits_last = PECross_51_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_67_multiply_io_input_io_actOut_ready = PECross_68_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_67_multiply_io_input_io_weiOut_ready = PECross_83_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_68_clock = clock;
  assign PECross_68_reset = rst;
  assign PECross_68_multiply_io_input_io_sumIn_valid = PECross_67_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_68_multiply_io_input_io_sumIn_bits_x_0 = PECross_67_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_68_multiply_io_input_io_sumIn_bits_last = PECross_67_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_68_multiply_io_input_io_sumOut_ready = PECross_69_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_68_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_68_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_68_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_68_multiply_io_input_io_actIn_valid = PECross_67_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_68_multiply_io_input_io_actIn_bits_x_0 = PECross_67_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_68_multiply_io_input_io_actIn_bits_last = PECross_67_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_68_multiply_io_input_io_weiIn_valid = PECross_52_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_68_multiply_io_input_io_weiIn_bits_x_0 = PECross_52_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_68_multiply_io_input_io_weiIn_bits_last = PECross_52_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_68_multiply_io_input_io_actOut_ready = PECross_69_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_68_multiply_io_input_io_weiOut_ready = PECross_84_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_69_clock = clock;
  assign PECross_69_reset = rst;
  assign PECross_69_multiply_io_input_io_sumIn_valid = PECross_68_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_69_multiply_io_input_io_sumIn_bits_x_0 = PECross_68_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_69_multiply_io_input_io_sumIn_bits_last = PECross_68_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_69_multiply_io_input_io_sumOut_ready = PECross_70_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_69_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_69_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_69_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_69_multiply_io_input_io_actIn_valid = PECross_68_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_69_multiply_io_input_io_actIn_bits_x_0 = PECross_68_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_69_multiply_io_input_io_actIn_bits_last = PECross_68_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_69_multiply_io_input_io_weiIn_valid = PECross_53_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_69_multiply_io_input_io_weiIn_bits_x_0 = PECross_53_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_69_multiply_io_input_io_weiIn_bits_last = PECross_53_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_69_multiply_io_input_io_actOut_ready = PECross_70_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_69_multiply_io_input_io_weiOut_ready = PECross_85_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_70_clock = clock;
  assign PECross_70_reset = rst;
  assign PECross_70_multiply_io_input_io_sumIn_valid = PECross_69_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_70_multiply_io_input_io_sumIn_bits_x_0 = PECross_69_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_70_multiply_io_input_io_sumIn_bits_last = PECross_69_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_70_multiply_io_input_io_sumOut_ready = PECross_71_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_70_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_70_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_70_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_70_multiply_io_input_io_actIn_valid = PECross_69_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_70_multiply_io_input_io_actIn_bits_x_0 = PECross_69_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_70_multiply_io_input_io_actIn_bits_last = PECross_69_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_70_multiply_io_input_io_weiIn_valid = PECross_54_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_70_multiply_io_input_io_weiIn_bits_x_0 = PECross_54_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_70_multiply_io_input_io_weiIn_bits_last = PECross_54_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_70_multiply_io_input_io_actOut_ready = PECross_71_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_70_multiply_io_input_io_weiOut_ready = PECross_86_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_71_clock = clock;
  assign PECross_71_reset = rst;
  assign PECross_71_multiply_io_input_io_sumIn_valid = PECross_70_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_71_multiply_io_input_io_sumIn_bits_x_0 = PECross_70_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_71_multiply_io_input_io_sumIn_bits_last = PECross_70_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_71_multiply_io_input_io_sumOut_ready = PECross_72_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_71_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_71_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_71_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_71_multiply_io_input_io_actIn_valid = PECross_70_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_71_multiply_io_input_io_actIn_bits_x_0 = PECross_70_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_71_multiply_io_input_io_actIn_bits_last = PECross_70_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_71_multiply_io_input_io_weiIn_valid = PECross_55_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_71_multiply_io_input_io_weiIn_bits_x_0 = PECross_55_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_71_multiply_io_input_io_weiIn_bits_last = PECross_55_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_71_multiply_io_input_io_actOut_ready = PECross_72_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_71_multiply_io_input_io_weiOut_ready = PECross_87_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_72_clock = clock;
  assign PECross_72_reset = rst;
  assign PECross_72_multiply_io_input_io_sumIn_valid = PECross_71_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_72_multiply_io_input_io_sumIn_bits_x_0 = PECross_71_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_72_multiply_io_input_io_sumIn_bits_last = PECross_71_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_72_multiply_io_input_io_sumOut_ready = PECross_73_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_72_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_72_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_72_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_72_multiply_io_input_io_actIn_valid = PECross_71_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_72_multiply_io_input_io_actIn_bits_x_0 = PECross_71_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_72_multiply_io_input_io_actIn_bits_last = PECross_71_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_72_multiply_io_input_io_weiIn_valid = PECross_56_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_72_multiply_io_input_io_weiIn_bits_x_0 = PECross_56_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_72_multiply_io_input_io_weiIn_bits_last = PECross_56_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_72_multiply_io_input_io_actOut_ready = PECross_73_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_72_multiply_io_input_io_weiOut_ready = PECross_88_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_73_clock = clock;
  assign PECross_73_reset = rst;
  assign PECross_73_multiply_io_input_io_sumIn_valid = PECross_72_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_73_multiply_io_input_io_sumIn_bits_x_0 = PECross_72_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_73_multiply_io_input_io_sumIn_bits_last = PECross_72_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_73_multiply_io_input_io_sumOut_ready = PECross_74_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_73_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_73_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_73_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_73_multiply_io_input_io_actIn_valid = PECross_72_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_73_multiply_io_input_io_actIn_bits_x_0 = PECross_72_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_73_multiply_io_input_io_actIn_bits_last = PECross_72_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_73_multiply_io_input_io_weiIn_valid = PECross_57_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_73_multiply_io_input_io_weiIn_bits_x_0 = PECross_57_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_73_multiply_io_input_io_weiIn_bits_last = PECross_57_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_73_multiply_io_input_io_actOut_ready = PECross_74_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_73_multiply_io_input_io_weiOut_ready = PECross_89_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_74_clock = clock;
  assign PECross_74_reset = rst;
  assign PECross_74_multiply_io_input_io_sumIn_valid = PECross_73_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_74_multiply_io_input_io_sumIn_bits_x_0 = PECross_73_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_74_multiply_io_input_io_sumIn_bits_last = PECross_73_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_74_multiply_io_input_io_sumOut_ready = PECross_75_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_74_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_74_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_74_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_74_multiply_io_input_io_actIn_valid = PECross_73_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_74_multiply_io_input_io_actIn_bits_x_0 = PECross_73_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_74_multiply_io_input_io_actIn_bits_last = PECross_73_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_74_multiply_io_input_io_weiIn_valid = PECross_58_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_74_multiply_io_input_io_weiIn_bits_x_0 = PECross_58_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_74_multiply_io_input_io_weiIn_bits_last = PECross_58_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_74_multiply_io_input_io_actOut_ready = PECross_75_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_74_multiply_io_input_io_weiOut_ready = PECross_90_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_75_clock = clock;
  assign PECross_75_reset = rst;
  assign PECross_75_multiply_io_input_io_sumIn_valid = PECross_74_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_75_multiply_io_input_io_sumIn_bits_x_0 = PECross_74_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_75_multiply_io_input_io_sumIn_bits_last = PECross_74_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_75_multiply_io_input_io_sumOut_ready = PECross_76_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_75_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_75_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_75_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_75_multiply_io_input_io_actIn_valid = PECross_74_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_75_multiply_io_input_io_actIn_bits_x_0 = PECross_74_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_75_multiply_io_input_io_actIn_bits_last = PECross_74_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_75_multiply_io_input_io_weiIn_valid = PECross_59_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_75_multiply_io_input_io_weiIn_bits_x_0 = PECross_59_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_75_multiply_io_input_io_weiIn_bits_last = PECross_59_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_75_multiply_io_input_io_actOut_ready = PECross_76_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_75_multiply_io_input_io_weiOut_ready = PECross_91_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_76_clock = clock;
  assign PECross_76_reset = rst;
  assign PECross_76_multiply_io_input_io_sumIn_valid = PECross_75_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_76_multiply_io_input_io_sumIn_bits_x_0 = PECross_75_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_76_multiply_io_input_io_sumIn_bits_last = PECross_75_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_76_multiply_io_input_io_sumOut_ready = PECross_77_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_76_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_76_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_76_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_76_multiply_io_input_io_actIn_valid = PECross_75_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_76_multiply_io_input_io_actIn_bits_x_0 = PECross_75_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_76_multiply_io_input_io_actIn_bits_last = PECross_75_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_76_multiply_io_input_io_weiIn_valid = PECross_60_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_76_multiply_io_input_io_weiIn_bits_x_0 = PECross_60_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_76_multiply_io_input_io_weiIn_bits_last = PECross_60_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_76_multiply_io_input_io_actOut_ready = PECross_77_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_76_multiply_io_input_io_weiOut_ready = PECross_92_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_77_clock = clock;
  assign PECross_77_reset = rst;
  assign PECross_77_multiply_io_input_io_sumIn_valid = PECross_76_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_77_multiply_io_input_io_sumIn_bits_x_0 = PECross_76_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_77_multiply_io_input_io_sumIn_bits_last = PECross_76_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_77_multiply_io_input_io_sumOut_ready = PECross_78_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_77_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_77_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_77_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_77_multiply_io_input_io_actIn_valid = PECross_76_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_77_multiply_io_input_io_actIn_bits_x_0 = PECross_76_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_77_multiply_io_input_io_actIn_bits_last = PECross_76_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_77_multiply_io_input_io_weiIn_valid = PECross_61_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_77_multiply_io_input_io_weiIn_bits_x_0 = PECross_61_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_77_multiply_io_input_io_weiIn_bits_last = PECross_61_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_77_multiply_io_input_io_actOut_ready = PECross_78_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_77_multiply_io_input_io_weiOut_ready = PECross_93_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_78_clock = clock;
  assign PECross_78_reset = rst;
  assign PECross_78_multiply_io_input_io_sumIn_valid = PECross_77_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_78_multiply_io_input_io_sumIn_bits_x_0 = PECross_77_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_78_multiply_io_input_io_sumIn_bits_last = PECross_77_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_78_multiply_io_input_io_sumOut_ready = PECross_79_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_78_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_78_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_78_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_78_multiply_io_input_io_actIn_valid = PECross_77_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_78_multiply_io_input_io_actIn_bits_x_0 = PECross_77_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_78_multiply_io_input_io_actIn_bits_last = PECross_77_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_78_multiply_io_input_io_weiIn_valid = PECross_62_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_78_multiply_io_input_io_weiIn_bits_x_0 = PECross_62_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_78_multiply_io_input_io_weiIn_bits_last = PECross_62_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_78_multiply_io_input_io_actOut_ready = PECross_79_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_78_multiply_io_input_io_weiOut_ready = PECross_94_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_79_clock = clock;
  assign PECross_79_reset = rst;
  assign PECross_79_multiply_io_input_io_sumIn_valid = PECross_78_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_79_multiply_io_input_io_sumIn_bits_x_0 = PECross_78_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_79_multiply_io_input_io_sumIn_bits_last = PECross_78_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_79_multiply_io_input_io_sumOut_ready = io_sumOut_4_ready; // @[mac.scala 45:29]
  assign PECross_79_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_79_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_79_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_79_multiply_io_input_io_actIn_valid = PECross_78_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_79_multiply_io_input_io_actIn_bits_x_0 = PECross_78_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_79_multiply_io_input_io_actIn_bits_last = PECross_78_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_79_multiply_io_input_io_weiIn_valid = PECross_63_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_79_multiply_io_input_io_weiIn_bits_x_0 = PECross_63_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_79_multiply_io_input_io_weiIn_bits_last = PECross_63_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_79_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_79_multiply_io_input_io_weiOut_ready = PECross_95_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_80_clock = clock;
  assign PECross_80_reset = rst;
  assign PECross_80_multiply_io_input_io_sumIn_valid = io_sumIn_5_valid; // @[mac.scala 33:28]
  assign PECross_80_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_5_bits_x_0; // @[mac.scala 33:28]
  assign PECross_80_multiply_io_input_io_sumIn_bits_last = io_sumIn_5_bits_last; // @[mac.scala 33:28]
  assign PECross_80_multiply_io_input_io_sumOut_ready = PECross_81_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_80_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_80_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_80_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_80_multiply_io_input_io_actIn_valid = io_actIn_5_valid; // @[mac.scala 32:28]
  assign PECross_80_multiply_io_input_io_actIn_bits_x_0 = io_actIn_5_bits_x_0; // @[mac.scala 32:28]
  assign PECross_80_multiply_io_input_io_actIn_bits_last = io_actIn_5_bits_last; // @[mac.scala 32:28]
  assign PECross_80_multiply_io_input_io_weiIn_valid = PECross_64_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_80_multiply_io_input_io_weiIn_bits_x_0 = PECross_64_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_80_multiply_io_input_io_weiIn_bits_last = PECross_64_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_80_multiply_io_input_io_actOut_ready = PECross_81_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_80_multiply_io_input_io_weiOut_ready = PECross_96_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_81_clock = clock;
  assign PECross_81_reset = rst;
  assign PECross_81_multiply_io_input_io_sumIn_valid = PECross_80_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_81_multiply_io_input_io_sumIn_bits_x_0 = PECross_80_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_81_multiply_io_input_io_sumIn_bits_last = PECross_80_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_81_multiply_io_input_io_sumOut_ready = PECross_82_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_81_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_81_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_81_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_81_multiply_io_input_io_actIn_valid = PECross_80_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_81_multiply_io_input_io_actIn_bits_x_0 = PECross_80_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_81_multiply_io_input_io_actIn_bits_last = PECross_80_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_81_multiply_io_input_io_weiIn_valid = PECross_65_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_81_multiply_io_input_io_weiIn_bits_x_0 = PECross_65_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_81_multiply_io_input_io_weiIn_bits_last = PECross_65_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_81_multiply_io_input_io_actOut_ready = PECross_82_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_81_multiply_io_input_io_weiOut_ready = PECross_97_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_82_clock = clock;
  assign PECross_82_reset = rst;
  assign PECross_82_multiply_io_input_io_sumIn_valid = PECross_81_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_82_multiply_io_input_io_sumIn_bits_x_0 = PECross_81_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_82_multiply_io_input_io_sumIn_bits_last = PECross_81_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_82_multiply_io_input_io_sumOut_ready = PECross_83_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_82_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_82_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_82_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_82_multiply_io_input_io_actIn_valid = PECross_81_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_82_multiply_io_input_io_actIn_bits_x_0 = PECross_81_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_82_multiply_io_input_io_actIn_bits_last = PECross_81_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_82_multiply_io_input_io_weiIn_valid = PECross_66_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_82_multiply_io_input_io_weiIn_bits_x_0 = PECross_66_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_82_multiply_io_input_io_weiIn_bits_last = PECross_66_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_82_multiply_io_input_io_actOut_ready = PECross_83_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_82_multiply_io_input_io_weiOut_ready = PECross_98_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_83_clock = clock;
  assign PECross_83_reset = rst;
  assign PECross_83_multiply_io_input_io_sumIn_valid = PECross_82_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_83_multiply_io_input_io_sumIn_bits_x_0 = PECross_82_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_83_multiply_io_input_io_sumIn_bits_last = PECross_82_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_83_multiply_io_input_io_sumOut_ready = PECross_84_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_83_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_83_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_83_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_83_multiply_io_input_io_actIn_valid = PECross_82_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_83_multiply_io_input_io_actIn_bits_x_0 = PECross_82_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_83_multiply_io_input_io_actIn_bits_last = PECross_82_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_83_multiply_io_input_io_weiIn_valid = PECross_67_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_83_multiply_io_input_io_weiIn_bits_x_0 = PECross_67_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_83_multiply_io_input_io_weiIn_bits_last = PECross_67_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_83_multiply_io_input_io_actOut_ready = PECross_84_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_83_multiply_io_input_io_weiOut_ready = PECross_99_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_84_clock = clock;
  assign PECross_84_reset = rst;
  assign PECross_84_multiply_io_input_io_sumIn_valid = PECross_83_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_84_multiply_io_input_io_sumIn_bits_x_0 = PECross_83_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_84_multiply_io_input_io_sumIn_bits_last = PECross_83_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_84_multiply_io_input_io_sumOut_ready = PECross_85_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_84_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_84_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_84_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_84_multiply_io_input_io_actIn_valid = PECross_83_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_84_multiply_io_input_io_actIn_bits_x_0 = PECross_83_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_84_multiply_io_input_io_actIn_bits_last = PECross_83_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_84_multiply_io_input_io_weiIn_valid = PECross_68_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_84_multiply_io_input_io_weiIn_bits_x_0 = PECross_68_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_84_multiply_io_input_io_weiIn_bits_last = PECross_68_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_84_multiply_io_input_io_actOut_ready = PECross_85_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_84_multiply_io_input_io_weiOut_ready = PECross_100_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_85_clock = clock;
  assign PECross_85_reset = rst;
  assign PECross_85_multiply_io_input_io_sumIn_valid = PECross_84_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_85_multiply_io_input_io_sumIn_bits_x_0 = PECross_84_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_85_multiply_io_input_io_sumIn_bits_last = PECross_84_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_85_multiply_io_input_io_sumOut_ready = PECross_86_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_85_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_85_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_85_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_85_multiply_io_input_io_actIn_valid = PECross_84_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_85_multiply_io_input_io_actIn_bits_x_0 = PECross_84_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_85_multiply_io_input_io_actIn_bits_last = PECross_84_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_85_multiply_io_input_io_weiIn_valid = PECross_69_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_85_multiply_io_input_io_weiIn_bits_x_0 = PECross_69_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_85_multiply_io_input_io_weiIn_bits_last = PECross_69_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_85_multiply_io_input_io_actOut_ready = PECross_86_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_85_multiply_io_input_io_weiOut_ready = PECross_101_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_86_clock = clock;
  assign PECross_86_reset = rst;
  assign PECross_86_multiply_io_input_io_sumIn_valid = PECross_85_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_86_multiply_io_input_io_sumIn_bits_x_0 = PECross_85_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_86_multiply_io_input_io_sumIn_bits_last = PECross_85_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_86_multiply_io_input_io_sumOut_ready = PECross_87_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_86_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_86_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_86_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_86_multiply_io_input_io_actIn_valid = PECross_85_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_86_multiply_io_input_io_actIn_bits_x_0 = PECross_85_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_86_multiply_io_input_io_actIn_bits_last = PECross_85_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_86_multiply_io_input_io_weiIn_valid = PECross_70_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_86_multiply_io_input_io_weiIn_bits_x_0 = PECross_70_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_86_multiply_io_input_io_weiIn_bits_last = PECross_70_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_86_multiply_io_input_io_actOut_ready = PECross_87_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_86_multiply_io_input_io_weiOut_ready = PECross_102_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_87_clock = clock;
  assign PECross_87_reset = rst;
  assign PECross_87_multiply_io_input_io_sumIn_valid = PECross_86_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_87_multiply_io_input_io_sumIn_bits_x_0 = PECross_86_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_87_multiply_io_input_io_sumIn_bits_last = PECross_86_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_87_multiply_io_input_io_sumOut_ready = PECross_88_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_87_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_87_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_87_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_87_multiply_io_input_io_actIn_valid = PECross_86_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_87_multiply_io_input_io_actIn_bits_x_0 = PECross_86_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_87_multiply_io_input_io_actIn_bits_last = PECross_86_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_87_multiply_io_input_io_weiIn_valid = PECross_71_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_87_multiply_io_input_io_weiIn_bits_x_0 = PECross_71_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_87_multiply_io_input_io_weiIn_bits_last = PECross_71_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_87_multiply_io_input_io_actOut_ready = PECross_88_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_87_multiply_io_input_io_weiOut_ready = PECross_103_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_88_clock = clock;
  assign PECross_88_reset = rst;
  assign PECross_88_multiply_io_input_io_sumIn_valid = PECross_87_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_88_multiply_io_input_io_sumIn_bits_x_0 = PECross_87_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_88_multiply_io_input_io_sumIn_bits_last = PECross_87_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_88_multiply_io_input_io_sumOut_ready = PECross_89_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_88_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_88_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_88_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_88_multiply_io_input_io_actIn_valid = PECross_87_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_88_multiply_io_input_io_actIn_bits_x_0 = PECross_87_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_88_multiply_io_input_io_actIn_bits_last = PECross_87_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_88_multiply_io_input_io_weiIn_valid = PECross_72_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_88_multiply_io_input_io_weiIn_bits_x_0 = PECross_72_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_88_multiply_io_input_io_weiIn_bits_last = PECross_72_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_88_multiply_io_input_io_actOut_ready = PECross_89_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_88_multiply_io_input_io_weiOut_ready = PECross_104_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_89_clock = clock;
  assign PECross_89_reset = rst;
  assign PECross_89_multiply_io_input_io_sumIn_valid = PECross_88_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_89_multiply_io_input_io_sumIn_bits_x_0 = PECross_88_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_89_multiply_io_input_io_sumIn_bits_last = PECross_88_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_89_multiply_io_input_io_sumOut_ready = PECross_90_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_89_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_89_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_89_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_89_multiply_io_input_io_actIn_valid = PECross_88_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_89_multiply_io_input_io_actIn_bits_x_0 = PECross_88_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_89_multiply_io_input_io_actIn_bits_last = PECross_88_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_89_multiply_io_input_io_weiIn_valid = PECross_73_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_89_multiply_io_input_io_weiIn_bits_x_0 = PECross_73_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_89_multiply_io_input_io_weiIn_bits_last = PECross_73_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_89_multiply_io_input_io_actOut_ready = PECross_90_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_89_multiply_io_input_io_weiOut_ready = PECross_105_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_90_clock = clock;
  assign PECross_90_reset = rst;
  assign PECross_90_multiply_io_input_io_sumIn_valid = PECross_89_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_90_multiply_io_input_io_sumIn_bits_x_0 = PECross_89_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_90_multiply_io_input_io_sumIn_bits_last = PECross_89_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_90_multiply_io_input_io_sumOut_ready = PECross_91_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_90_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_90_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_90_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_90_multiply_io_input_io_actIn_valid = PECross_89_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_90_multiply_io_input_io_actIn_bits_x_0 = PECross_89_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_90_multiply_io_input_io_actIn_bits_last = PECross_89_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_90_multiply_io_input_io_weiIn_valid = PECross_74_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_90_multiply_io_input_io_weiIn_bits_x_0 = PECross_74_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_90_multiply_io_input_io_weiIn_bits_last = PECross_74_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_90_multiply_io_input_io_actOut_ready = PECross_91_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_90_multiply_io_input_io_weiOut_ready = PECross_106_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_91_clock = clock;
  assign PECross_91_reset = rst;
  assign PECross_91_multiply_io_input_io_sumIn_valid = PECross_90_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_91_multiply_io_input_io_sumIn_bits_x_0 = PECross_90_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_91_multiply_io_input_io_sumIn_bits_last = PECross_90_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_91_multiply_io_input_io_sumOut_ready = PECross_92_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_91_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_91_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_91_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_91_multiply_io_input_io_actIn_valid = PECross_90_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_91_multiply_io_input_io_actIn_bits_x_0 = PECross_90_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_91_multiply_io_input_io_actIn_bits_last = PECross_90_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_91_multiply_io_input_io_weiIn_valid = PECross_75_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_91_multiply_io_input_io_weiIn_bits_x_0 = PECross_75_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_91_multiply_io_input_io_weiIn_bits_last = PECross_75_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_91_multiply_io_input_io_actOut_ready = PECross_92_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_91_multiply_io_input_io_weiOut_ready = PECross_107_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_92_clock = clock;
  assign PECross_92_reset = rst;
  assign PECross_92_multiply_io_input_io_sumIn_valid = PECross_91_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_92_multiply_io_input_io_sumIn_bits_x_0 = PECross_91_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_92_multiply_io_input_io_sumIn_bits_last = PECross_91_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_92_multiply_io_input_io_sumOut_ready = PECross_93_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_92_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_92_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_92_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_92_multiply_io_input_io_actIn_valid = PECross_91_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_92_multiply_io_input_io_actIn_bits_x_0 = PECross_91_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_92_multiply_io_input_io_actIn_bits_last = PECross_91_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_92_multiply_io_input_io_weiIn_valid = PECross_76_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_92_multiply_io_input_io_weiIn_bits_x_0 = PECross_76_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_92_multiply_io_input_io_weiIn_bits_last = PECross_76_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_92_multiply_io_input_io_actOut_ready = PECross_93_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_92_multiply_io_input_io_weiOut_ready = PECross_108_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_93_clock = clock;
  assign PECross_93_reset = rst;
  assign PECross_93_multiply_io_input_io_sumIn_valid = PECross_92_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_93_multiply_io_input_io_sumIn_bits_x_0 = PECross_92_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_93_multiply_io_input_io_sumIn_bits_last = PECross_92_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_93_multiply_io_input_io_sumOut_ready = PECross_94_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_93_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_93_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_93_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_93_multiply_io_input_io_actIn_valid = PECross_92_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_93_multiply_io_input_io_actIn_bits_x_0 = PECross_92_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_93_multiply_io_input_io_actIn_bits_last = PECross_92_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_93_multiply_io_input_io_weiIn_valid = PECross_77_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_93_multiply_io_input_io_weiIn_bits_x_0 = PECross_77_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_93_multiply_io_input_io_weiIn_bits_last = PECross_77_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_93_multiply_io_input_io_actOut_ready = PECross_94_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_93_multiply_io_input_io_weiOut_ready = PECross_109_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_94_clock = clock;
  assign PECross_94_reset = rst;
  assign PECross_94_multiply_io_input_io_sumIn_valid = PECross_93_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_94_multiply_io_input_io_sumIn_bits_x_0 = PECross_93_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_94_multiply_io_input_io_sumIn_bits_last = PECross_93_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_94_multiply_io_input_io_sumOut_ready = PECross_95_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_94_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_94_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_94_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_94_multiply_io_input_io_actIn_valid = PECross_93_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_94_multiply_io_input_io_actIn_bits_x_0 = PECross_93_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_94_multiply_io_input_io_actIn_bits_last = PECross_93_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_94_multiply_io_input_io_weiIn_valid = PECross_78_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_94_multiply_io_input_io_weiIn_bits_x_0 = PECross_78_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_94_multiply_io_input_io_weiIn_bits_last = PECross_78_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_94_multiply_io_input_io_actOut_ready = PECross_95_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_94_multiply_io_input_io_weiOut_ready = PECross_110_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_95_clock = clock;
  assign PECross_95_reset = rst;
  assign PECross_95_multiply_io_input_io_sumIn_valid = PECross_94_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_95_multiply_io_input_io_sumIn_bits_x_0 = PECross_94_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_95_multiply_io_input_io_sumIn_bits_last = PECross_94_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_95_multiply_io_input_io_sumOut_ready = io_sumOut_5_ready; // @[mac.scala 45:29]
  assign PECross_95_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_95_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_95_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_95_multiply_io_input_io_actIn_valid = PECross_94_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_95_multiply_io_input_io_actIn_bits_x_0 = PECross_94_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_95_multiply_io_input_io_actIn_bits_last = PECross_94_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_95_multiply_io_input_io_weiIn_valid = PECross_79_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_95_multiply_io_input_io_weiIn_bits_x_0 = PECross_79_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_95_multiply_io_input_io_weiIn_bits_last = PECross_79_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_95_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_95_multiply_io_input_io_weiOut_ready = PECross_111_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_96_clock = clock;
  assign PECross_96_reset = rst;
  assign PECross_96_multiply_io_input_io_sumIn_valid = io_sumIn_6_valid; // @[mac.scala 33:28]
  assign PECross_96_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_6_bits_x_0; // @[mac.scala 33:28]
  assign PECross_96_multiply_io_input_io_sumIn_bits_last = io_sumIn_6_bits_last; // @[mac.scala 33:28]
  assign PECross_96_multiply_io_input_io_sumOut_ready = PECross_97_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_96_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_96_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_96_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_96_multiply_io_input_io_actIn_valid = io_actIn_6_valid; // @[mac.scala 32:28]
  assign PECross_96_multiply_io_input_io_actIn_bits_x_0 = io_actIn_6_bits_x_0; // @[mac.scala 32:28]
  assign PECross_96_multiply_io_input_io_actIn_bits_last = io_actIn_6_bits_last; // @[mac.scala 32:28]
  assign PECross_96_multiply_io_input_io_weiIn_valid = PECross_80_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_96_multiply_io_input_io_weiIn_bits_x_0 = PECross_80_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_96_multiply_io_input_io_weiIn_bits_last = PECross_80_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_96_multiply_io_input_io_actOut_ready = PECross_97_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_96_multiply_io_input_io_weiOut_ready = PECross_112_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_97_clock = clock;
  assign PECross_97_reset = rst;
  assign PECross_97_multiply_io_input_io_sumIn_valid = PECross_96_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_97_multiply_io_input_io_sumIn_bits_x_0 = PECross_96_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_97_multiply_io_input_io_sumIn_bits_last = PECross_96_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_97_multiply_io_input_io_sumOut_ready = PECross_98_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_97_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_97_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_97_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_97_multiply_io_input_io_actIn_valid = PECross_96_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_97_multiply_io_input_io_actIn_bits_x_0 = PECross_96_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_97_multiply_io_input_io_actIn_bits_last = PECross_96_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_97_multiply_io_input_io_weiIn_valid = PECross_81_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_97_multiply_io_input_io_weiIn_bits_x_0 = PECross_81_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_97_multiply_io_input_io_weiIn_bits_last = PECross_81_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_97_multiply_io_input_io_actOut_ready = PECross_98_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_97_multiply_io_input_io_weiOut_ready = PECross_113_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_98_clock = clock;
  assign PECross_98_reset = rst;
  assign PECross_98_multiply_io_input_io_sumIn_valid = PECross_97_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_98_multiply_io_input_io_sumIn_bits_x_0 = PECross_97_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_98_multiply_io_input_io_sumIn_bits_last = PECross_97_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_98_multiply_io_input_io_sumOut_ready = PECross_99_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_98_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_98_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_98_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_98_multiply_io_input_io_actIn_valid = PECross_97_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_98_multiply_io_input_io_actIn_bits_x_0 = PECross_97_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_98_multiply_io_input_io_actIn_bits_last = PECross_97_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_98_multiply_io_input_io_weiIn_valid = PECross_82_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_98_multiply_io_input_io_weiIn_bits_x_0 = PECross_82_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_98_multiply_io_input_io_weiIn_bits_last = PECross_82_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_98_multiply_io_input_io_actOut_ready = PECross_99_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_98_multiply_io_input_io_weiOut_ready = PECross_114_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_99_clock = clock;
  assign PECross_99_reset = rst;
  assign PECross_99_multiply_io_input_io_sumIn_valid = PECross_98_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_99_multiply_io_input_io_sumIn_bits_x_0 = PECross_98_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_99_multiply_io_input_io_sumIn_bits_last = PECross_98_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_99_multiply_io_input_io_sumOut_ready = PECross_100_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_99_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_99_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_99_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_99_multiply_io_input_io_actIn_valid = PECross_98_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_99_multiply_io_input_io_actIn_bits_x_0 = PECross_98_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_99_multiply_io_input_io_actIn_bits_last = PECross_98_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_99_multiply_io_input_io_weiIn_valid = PECross_83_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_99_multiply_io_input_io_weiIn_bits_x_0 = PECross_83_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_99_multiply_io_input_io_weiIn_bits_last = PECross_83_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_99_multiply_io_input_io_actOut_ready = PECross_100_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_99_multiply_io_input_io_weiOut_ready = PECross_115_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_100_clock = clock;
  assign PECross_100_reset = rst;
  assign PECross_100_multiply_io_input_io_sumIn_valid = PECross_99_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_100_multiply_io_input_io_sumIn_bits_x_0 = PECross_99_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_100_multiply_io_input_io_sumIn_bits_last = PECross_99_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_100_multiply_io_input_io_sumOut_ready = PECross_101_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_100_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_100_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_100_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_100_multiply_io_input_io_actIn_valid = PECross_99_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_100_multiply_io_input_io_actIn_bits_x_0 = PECross_99_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_100_multiply_io_input_io_actIn_bits_last = PECross_99_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_100_multiply_io_input_io_weiIn_valid = PECross_84_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_100_multiply_io_input_io_weiIn_bits_x_0 = PECross_84_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_100_multiply_io_input_io_weiIn_bits_last = PECross_84_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_100_multiply_io_input_io_actOut_ready = PECross_101_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_100_multiply_io_input_io_weiOut_ready = PECross_116_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_101_clock = clock;
  assign PECross_101_reset = rst;
  assign PECross_101_multiply_io_input_io_sumIn_valid = PECross_100_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_101_multiply_io_input_io_sumIn_bits_x_0 = PECross_100_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_101_multiply_io_input_io_sumIn_bits_last = PECross_100_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_101_multiply_io_input_io_sumOut_ready = PECross_102_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_101_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_101_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_101_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_101_multiply_io_input_io_actIn_valid = PECross_100_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_101_multiply_io_input_io_actIn_bits_x_0 = PECross_100_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_101_multiply_io_input_io_actIn_bits_last = PECross_100_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_101_multiply_io_input_io_weiIn_valid = PECross_85_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_101_multiply_io_input_io_weiIn_bits_x_0 = PECross_85_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_101_multiply_io_input_io_weiIn_bits_last = PECross_85_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_101_multiply_io_input_io_actOut_ready = PECross_102_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_101_multiply_io_input_io_weiOut_ready = PECross_117_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_102_clock = clock;
  assign PECross_102_reset = rst;
  assign PECross_102_multiply_io_input_io_sumIn_valid = PECross_101_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_102_multiply_io_input_io_sumIn_bits_x_0 = PECross_101_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_102_multiply_io_input_io_sumIn_bits_last = PECross_101_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_102_multiply_io_input_io_sumOut_ready = PECross_103_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_102_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_102_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_102_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_102_multiply_io_input_io_actIn_valid = PECross_101_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_102_multiply_io_input_io_actIn_bits_x_0 = PECross_101_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_102_multiply_io_input_io_actIn_bits_last = PECross_101_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_102_multiply_io_input_io_weiIn_valid = PECross_86_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_102_multiply_io_input_io_weiIn_bits_x_0 = PECross_86_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_102_multiply_io_input_io_weiIn_bits_last = PECross_86_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_102_multiply_io_input_io_actOut_ready = PECross_103_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_102_multiply_io_input_io_weiOut_ready = PECross_118_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_103_clock = clock;
  assign PECross_103_reset = rst;
  assign PECross_103_multiply_io_input_io_sumIn_valid = PECross_102_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_103_multiply_io_input_io_sumIn_bits_x_0 = PECross_102_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_103_multiply_io_input_io_sumIn_bits_last = PECross_102_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_103_multiply_io_input_io_sumOut_ready = PECross_104_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_103_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_103_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_103_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_103_multiply_io_input_io_actIn_valid = PECross_102_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_103_multiply_io_input_io_actIn_bits_x_0 = PECross_102_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_103_multiply_io_input_io_actIn_bits_last = PECross_102_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_103_multiply_io_input_io_weiIn_valid = PECross_87_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_103_multiply_io_input_io_weiIn_bits_x_0 = PECross_87_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_103_multiply_io_input_io_weiIn_bits_last = PECross_87_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_103_multiply_io_input_io_actOut_ready = PECross_104_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_103_multiply_io_input_io_weiOut_ready = PECross_119_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_104_clock = clock;
  assign PECross_104_reset = rst;
  assign PECross_104_multiply_io_input_io_sumIn_valid = PECross_103_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_104_multiply_io_input_io_sumIn_bits_x_0 = PECross_103_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_104_multiply_io_input_io_sumIn_bits_last = PECross_103_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_104_multiply_io_input_io_sumOut_ready = PECross_105_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_104_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_104_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_104_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_104_multiply_io_input_io_actIn_valid = PECross_103_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_104_multiply_io_input_io_actIn_bits_x_0 = PECross_103_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_104_multiply_io_input_io_actIn_bits_last = PECross_103_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_104_multiply_io_input_io_weiIn_valid = PECross_88_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_104_multiply_io_input_io_weiIn_bits_x_0 = PECross_88_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_104_multiply_io_input_io_weiIn_bits_last = PECross_88_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_104_multiply_io_input_io_actOut_ready = PECross_105_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_104_multiply_io_input_io_weiOut_ready = PECross_120_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_105_clock = clock;
  assign PECross_105_reset = rst;
  assign PECross_105_multiply_io_input_io_sumIn_valid = PECross_104_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_105_multiply_io_input_io_sumIn_bits_x_0 = PECross_104_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_105_multiply_io_input_io_sumIn_bits_last = PECross_104_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_105_multiply_io_input_io_sumOut_ready = PECross_106_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_105_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_105_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_105_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_105_multiply_io_input_io_actIn_valid = PECross_104_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_105_multiply_io_input_io_actIn_bits_x_0 = PECross_104_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_105_multiply_io_input_io_actIn_bits_last = PECross_104_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_105_multiply_io_input_io_weiIn_valid = PECross_89_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_105_multiply_io_input_io_weiIn_bits_x_0 = PECross_89_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_105_multiply_io_input_io_weiIn_bits_last = PECross_89_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_105_multiply_io_input_io_actOut_ready = PECross_106_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_105_multiply_io_input_io_weiOut_ready = PECross_121_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_106_clock = clock;
  assign PECross_106_reset = rst;
  assign PECross_106_multiply_io_input_io_sumIn_valid = PECross_105_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_106_multiply_io_input_io_sumIn_bits_x_0 = PECross_105_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_106_multiply_io_input_io_sumIn_bits_last = PECross_105_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_106_multiply_io_input_io_sumOut_ready = PECross_107_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_106_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_106_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_106_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_106_multiply_io_input_io_actIn_valid = PECross_105_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_106_multiply_io_input_io_actIn_bits_x_0 = PECross_105_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_106_multiply_io_input_io_actIn_bits_last = PECross_105_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_106_multiply_io_input_io_weiIn_valid = PECross_90_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_106_multiply_io_input_io_weiIn_bits_x_0 = PECross_90_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_106_multiply_io_input_io_weiIn_bits_last = PECross_90_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_106_multiply_io_input_io_actOut_ready = PECross_107_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_106_multiply_io_input_io_weiOut_ready = PECross_122_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_107_clock = clock;
  assign PECross_107_reset = rst;
  assign PECross_107_multiply_io_input_io_sumIn_valid = PECross_106_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_107_multiply_io_input_io_sumIn_bits_x_0 = PECross_106_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_107_multiply_io_input_io_sumIn_bits_last = PECross_106_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_107_multiply_io_input_io_sumOut_ready = PECross_108_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_107_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_107_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_107_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_107_multiply_io_input_io_actIn_valid = PECross_106_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_107_multiply_io_input_io_actIn_bits_x_0 = PECross_106_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_107_multiply_io_input_io_actIn_bits_last = PECross_106_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_107_multiply_io_input_io_weiIn_valid = PECross_91_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_107_multiply_io_input_io_weiIn_bits_x_0 = PECross_91_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_107_multiply_io_input_io_weiIn_bits_last = PECross_91_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_107_multiply_io_input_io_actOut_ready = PECross_108_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_107_multiply_io_input_io_weiOut_ready = PECross_123_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_108_clock = clock;
  assign PECross_108_reset = rst;
  assign PECross_108_multiply_io_input_io_sumIn_valid = PECross_107_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_108_multiply_io_input_io_sumIn_bits_x_0 = PECross_107_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_108_multiply_io_input_io_sumIn_bits_last = PECross_107_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_108_multiply_io_input_io_sumOut_ready = PECross_109_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_108_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_108_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_108_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_108_multiply_io_input_io_actIn_valid = PECross_107_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_108_multiply_io_input_io_actIn_bits_x_0 = PECross_107_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_108_multiply_io_input_io_actIn_bits_last = PECross_107_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_108_multiply_io_input_io_weiIn_valid = PECross_92_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_108_multiply_io_input_io_weiIn_bits_x_0 = PECross_92_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_108_multiply_io_input_io_weiIn_bits_last = PECross_92_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_108_multiply_io_input_io_actOut_ready = PECross_109_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_108_multiply_io_input_io_weiOut_ready = PECross_124_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_109_clock = clock;
  assign PECross_109_reset = rst;
  assign PECross_109_multiply_io_input_io_sumIn_valid = PECross_108_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_109_multiply_io_input_io_sumIn_bits_x_0 = PECross_108_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_109_multiply_io_input_io_sumIn_bits_last = PECross_108_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_109_multiply_io_input_io_sumOut_ready = PECross_110_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_109_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_109_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_109_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_109_multiply_io_input_io_actIn_valid = PECross_108_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_109_multiply_io_input_io_actIn_bits_x_0 = PECross_108_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_109_multiply_io_input_io_actIn_bits_last = PECross_108_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_109_multiply_io_input_io_weiIn_valid = PECross_93_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_109_multiply_io_input_io_weiIn_bits_x_0 = PECross_93_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_109_multiply_io_input_io_weiIn_bits_last = PECross_93_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_109_multiply_io_input_io_actOut_ready = PECross_110_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_109_multiply_io_input_io_weiOut_ready = PECross_125_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_110_clock = clock;
  assign PECross_110_reset = rst;
  assign PECross_110_multiply_io_input_io_sumIn_valid = PECross_109_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_110_multiply_io_input_io_sumIn_bits_x_0 = PECross_109_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_110_multiply_io_input_io_sumIn_bits_last = PECross_109_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_110_multiply_io_input_io_sumOut_ready = PECross_111_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_110_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_110_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_110_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_110_multiply_io_input_io_actIn_valid = PECross_109_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_110_multiply_io_input_io_actIn_bits_x_0 = PECross_109_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_110_multiply_io_input_io_actIn_bits_last = PECross_109_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_110_multiply_io_input_io_weiIn_valid = PECross_94_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_110_multiply_io_input_io_weiIn_bits_x_0 = PECross_94_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_110_multiply_io_input_io_weiIn_bits_last = PECross_94_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_110_multiply_io_input_io_actOut_ready = PECross_111_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_110_multiply_io_input_io_weiOut_ready = PECross_126_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_111_clock = clock;
  assign PECross_111_reset = rst;
  assign PECross_111_multiply_io_input_io_sumIn_valid = PECross_110_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_111_multiply_io_input_io_sumIn_bits_x_0 = PECross_110_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_111_multiply_io_input_io_sumIn_bits_last = PECross_110_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_111_multiply_io_input_io_sumOut_ready = io_sumOut_6_ready; // @[mac.scala 45:29]
  assign PECross_111_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_111_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_111_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_111_multiply_io_input_io_actIn_valid = PECross_110_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_111_multiply_io_input_io_actIn_bits_x_0 = PECross_110_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_111_multiply_io_input_io_actIn_bits_last = PECross_110_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_111_multiply_io_input_io_weiIn_valid = PECross_95_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_111_multiply_io_input_io_weiIn_bits_x_0 = PECross_95_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_111_multiply_io_input_io_weiIn_bits_last = PECross_95_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_111_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_111_multiply_io_input_io_weiOut_ready = PECross_127_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_112_clock = clock;
  assign PECross_112_reset = rst;
  assign PECross_112_multiply_io_input_io_sumIn_valid = io_sumIn_7_valid; // @[mac.scala 33:28]
  assign PECross_112_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_7_bits_x_0; // @[mac.scala 33:28]
  assign PECross_112_multiply_io_input_io_sumIn_bits_last = io_sumIn_7_bits_last; // @[mac.scala 33:28]
  assign PECross_112_multiply_io_input_io_sumOut_ready = PECross_113_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_112_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_112_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_112_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_112_multiply_io_input_io_actIn_valid = io_actIn_7_valid; // @[mac.scala 32:28]
  assign PECross_112_multiply_io_input_io_actIn_bits_x_0 = io_actIn_7_bits_x_0; // @[mac.scala 32:28]
  assign PECross_112_multiply_io_input_io_actIn_bits_last = io_actIn_7_bits_last; // @[mac.scala 32:28]
  assign PECross_112_multiply_io_input_io_weiIn_valid = PECross_96_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_112_multiply_io_input_io_weiIn_bits_x_0 = PECross_96_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_112_multiply_io_input_io_weiIn_bits_last = PECross_96_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_112_multiply_io_input_io_actOut_ready = PECross_113_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_112_multiply_io_input_io_weiOut_ready = PECross_128_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_113_clock = clock;
  assign PECross_113_reset = rst;
  assign PECross_113_multiply_io_input_io_sumIn_valid = PECross_112_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_113_multiply_io_input_io_sumIn_bits_x_0 = PECross_112_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_113_multiply_io_input_io_sumIn_bits_last = PECross_112_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_113_multiply_io_input_io_sumOut_ready = PECross_114_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_113_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_113_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_113_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_113_multiply_io_input_io_actIn_valid = PECross_112_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_113_multiply_io_input_io_actIn_bits_x_0 = PECross_112_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_113_multiply_io_input_io_actIn_bits_last = PECross_112_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_113_multiply_io_input_io_weiIn_valid = PECross_97_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_113_multiply_io_input_io_weiIn_bits_x_0 = PECross_97_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_113_multiply_io_input_io_weiIn_bits_last = PECross_97_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_113_multiply_io_input_io_actOut_ready = PECross_114_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_113_multiply_io_input_io_weiOut_ready = PECross_129_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_114_clock = clock;
  assign PECross_114_reset = rst;
  assign PECross_114_multiply_io_input_io_sumIn_valid = PECross_113_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_114_multiply_io_input_io_sumIn_bits_x_0 = PECross_113_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_114_multiply_io_input_io_sumIn_bits_last = PECross_113_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_114_multiply_io_input_io_sumOut_ready = PECross_115_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_114_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_114_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_114_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_114_multiply_io_input_io_actIn_valid = PECross_113_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_114_multiply_io_input_io_actIn_bits_x_0 = PECross_113_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_114_multiply_io_input_io_actIn_bits_last = PECross_113_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_114_multiply_io_input_io_weiIn_valid = PECross_98_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_114_multiply_io_input_io_weiIn_bits_x_0 = PECross_98_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_114_multiply_io_input_io_weiIn_bits_last = PECross_98_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_114_multiply_io_input_io_actOut_ready = PECross_115_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_114_multiply_io_input_io_weiOut_ready = PECross_130_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_115_clock = clock;
  assign PECross_115_reset = rst;
  assign PECross_115_multiply_io_input_io_sumIn_valid = PECross_114_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_115_multiply_io_input_io_sumIn_bits_x_0 = PECross_114_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_115_multiply_io_input_io_sumIn_bits_last = PECross_114_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_115_multiply_io_input_io_sumOut_ready = PECross_116_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_115_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_115_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_115_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_115_multiply_io_input_io_actIn_valid = PECross_114_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_115_multiply_io_input_io_actIn_bits_x_0 = PECross_114_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_115_multiply_io_input_io_actIn_bits_last = PECross_114_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_115_multiply_io_input_io_weiIn_valid = PECross_99_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_115_multiply_io_input_io_weiIn_bits_x_0 = PECross_99_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_115_multiply_io_input_io_weiIn_bits_last = PECross_99_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_115_multiply_io_input_io_actOut_ready = PECross_116_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_115_multiply_io_input_io_weiOut_ready = PECross_131_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_116_clock = clock;
  assign PECross_116_reset = rst;
  assign PECross_116_multiply_io_input_io_sumIn_valid = PECross_115_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_116_multiply_io_input_io_sumIn_bits_x_0 = PECross_115_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_116_multiply_io_input_io_sumIn_bits_last = PECross_115_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_116_multiply_io_input_io_sumOut_ready = PECross_117_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_116_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_116_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_116_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_116_multiply_io_input_io_actIn_valid = PECross_115_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_116_multiply_io_input_io_actIn_bits_x_0 = PECross_115_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_116_multiply_io_input_io_actIn_bits_last = PECross_115_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_116_multiply_io_input_io_weiIn_valid = PECross_100_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_116_multiply_io_input_io_weiIn_bits_x_0 = PECross_100_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_116_multiply_io_input_io_weiIn_bits_last = PECross_100_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_116_multiply_io_input_io_actOut_ready = PECross_117_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_116_multiply_io_input_io_weiOut_ready = PECross_132_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_117_clock = clock;
  assign PECross_117_reset = rst;
  assign PECross_117_multiply_io_input_io_sumIn_valid = PECross_116_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_117_multiply_io_input_io_sumIn_bits_x_0 = PECross_116_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_117_multiply_io_input_io_sumIn_bits_last = PECross_116_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_117_multiply_io_input_io_sumOut_ready = PECross_118_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_117_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_117_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_117_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_117_multiply_io_input_io_actIn_valid = PECross_116_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_117_multiply_io_input_io_actIn_bits_x_0 = PECross_116_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_117_multiply_io_input_io_actIn_bits_last = PECross_116_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_117_multiply_io_input_io_weiIn_valid = PECross_101_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_117_multiply_io_input_io_weiIn_bits_x_0 = PECross_101_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_117_multiply_io_input_io_weiIn_bits_last = PECross_101_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_117_multiply_io_input_io_actOut_ready = PECross_118_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_117_multiply_io_input_io_weiOut_ready = PECross_133_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_118_clock = clock;
  assign PECross_118_reset = rst;
  assign PECross_118_multiply_io_input_io_sumIn_valid = PECross_117_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_118_multiply_io_input_io_sumIn_bits_x_0 = PECross_117_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_118_multiply_io_input_io_sumIn_bits_last = PECross_117_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_118_multiply_io_input_io_sumOut_ready = PECross_119_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_118_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_118_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_118_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_118_multiply_io_input_io_actIn_valid = PECross_117_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_118_multiply_io_input_io_actIn_bits_x_0 = PECross_117_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_118_multiply_io_input_io_actIn_bits_last = PECross_117_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_118_multiply_io_input_io_weiIn_valid = PECross_102_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_118_multiply_io_input_io_weiIn_bits_x_0 = PECross_102_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_118_multiply_io_input_io_weiIn_bits_last = PECross_102_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_118_multiply_io_input_io_actOut_ready = PECross_119_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_118_multiply_io_input_io_weiOut_ready = PECross_134_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_119_clock = clock;
  assign PECross_119_reset = rst;
  assign PECross_119_multiply_io_input_io_sumIn_valid = PECross_118_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_119_multiply_io_input_io_sumIn_bits_x_0 = PECross_118_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_119_multiply_io_input_io_sumIn_bits_last = PECross_118_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_119_multiply_io_input_io_sumOut_ready = PECross_120_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_119_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_119_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_119_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_119_multiply_io_input_io_actIn_valid = PECross_118_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_119_multiply_io_input_io_actIn_bits_x_0 = PECross_118_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_119_multiply_io_input_io_actIn_bits_last = PECross_118_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_119_multiply_io_input_io_weiIn_valid = PECross_103_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_119_multiply_io_input_io_weiIn_bits_x_0 = PECross_103_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_119_multiply_io_input_io_weiIn_bits_last = PECross_103_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_119_multiply_io_input_io_actOut_ready = PECross_120_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_119_multiply_io_input_io_weiOut_ready = PECross_135_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_120_clock = clock;
  assign PECross_120_reset = rst;
  assign PECross_120_multiply_io_input_io_sumIn_valid = PECross_119_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_120_multiply_io_input_io_sumIn_bits_x_0 = PECross_119_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_120_multiply_io_input_io_sumIn_bits_last = PECross_119_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_120_multiply_io_input_io_sumOut_ready = PECross_121_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_120_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_120_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_120_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_120_multiply_io_input_io_actIn_valid = PECross_119_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_120_multiply_io_input_io_actIn_bits_x_0 = PECross_119_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_120_multiply_io_input_io_actIn_bits_last = PECross_119_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_120_multiply_io_input_io_weiIn_valid = PECross_104_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_120_multiply_io_input_io_weiIn_bits_x_0 = PECross_104_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_120_multiply_io_input_io_weiIn_bits_last = PECross_104_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_120_multiply_io_input_io_actOut_ready = PECross_121_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_120_multiply_io_input_io_weiOut_ready = PECross_136_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_121_clock = clock;
  assign PECross_121_reset = rst;
  assign PECross_121_multiply_io_input_io_sumIn_valid = PECross_120_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_121_multiply_io_input_io_sumIn_bits_x_0 = PECross_120_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_121_multiply_io_input_io_sumIn_bits_last = PECross_120_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_121_multiply_io_input_io_sumOut_ready = PECross_122_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_121_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_121_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_121_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_121_multiply_io_input_io_actIn_valid = PECross_120_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_121_multiply_io_input_io_actIn_bits_x_0 = PECross_120_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_121_multiply_io_input_io_actIn_bits_last = PECross_120_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_121_multiply_io_input_io_weiIn_valid = PECross_105_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_121_multiply_io_input_io_weiIn_bits_x_0 = PECross_105_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_121_multiply_io_input_io_weiIn_bits_last = PECross_105_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_121_multiply_io_input_io_actOut_ready = PECross_122_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_121_multiply_io_input_io_weiOut_ready = PECross_137_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_122_clock = clock;
  assign PECross_122_reset = rst;
  assign PECross_122_multiply_io_input_io_sumIn_valid = PECross_121_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_122_multiply_io_input_io_sumIn_bits_x_0 = PECross_121_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_122_multiply_io_input_io_sumIn_bits_last = PECross_121_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_122_multiply_io_input_io_sumOut_ready = PECross_123_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_122_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_122_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_122_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_122_multiply_io_input_io_actIn_valid = PECross_121_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_122_multiply_io_input_io_actIn_bits_x_0 = PECross_121_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_122_multiply_io_input_io_actIn_bits_last = PECross_121_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_122_multiply_io_input_io_weiIn_valid = PECross_106_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_122_multiply_io_input_io_weiIn_bits_x_0 = PECross_106_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_122_multiply_io_input_io_weiIn_bits_last = PECross_106_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_122_multiply_io_input_io_actOut_ready = PECross_123_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_122_multiply_io_input_io_weiOut_ready = PECross_138_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_123_clock = clock;
  assign PECross_123_reset = rst;
  assign PECross_123_multiply_io_input_io_sumIn_valid = PECross_122_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_123_multiply_io_input_io_sumIn_bits_x_0 = PECross_122_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_123_multiply_io_input_io_sumIn_bits_last = PECross_122_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_123_multiply_io_input_io_sumOut_ready = PECross_124_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_123_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_123_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_123_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_123_multiply_io_input_io_actIn_valid = PECross_122_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_123_multiply_io_input_io_actIn_bits_x_0 = PECross_122_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_123_multiply_io_input_io_actIn_bits_last = PECross_122_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_123_multiply_io_input_io_weiIn_valid = PECross_107_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_123_multiply_io_input_io_weiIn_bits_x_0 = PECross_107_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_123_multiply_io_input_io_weiIn_bits_last = PECross_107_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_123_multiply_io_input_io_actOut_ready = PECross_124_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_123_multiply_io_input_io_weiOut_ready = PECross_139_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_124_clock = clock;
  assign PECross_124_reset = rst;
  assign PECross_124_multiply_io_input_io_sumIn_valid = PECross_123_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_124_multiply_io_input_io_sumIn_bits_x_0 = PECross_123_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_124_multiply_io_input_io_sumIn_bits_last = PECross_123_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_124_multiply_io_input_io_sumOut_ready = PECross_125_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_124_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_124_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_124_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_124_multiply_io_input_io_actIn_valid = PECross_123_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_124_multiply_io_input_io_actIn_bits_x_0 = PECross_123_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_124_multiply_io_input_io_actIn_bits_last = PECross_123_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_124_multiply_io_input_io_weiIn_valid = PECross_108_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_124_multiply_io_input_io_weiIn_bits_x_0 = PECross_108_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_124_multiply_io_input_io_weiIn_bits_last = PECross_108_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_124_multiply_io_input_io_actOut_ready = PECross_125_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_124_multiply_io_input_io_weiOut_ready = PECross_140_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_125_clock = clock;
  assign PECross_125_reset = rst;
  assign PECross_125_multiply_io_input_io_sumIn_valid = PECross_124_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_125_multiply_io_input_io_sumIn_bits_x_0 = PECross_124_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_125_multiply_io_input_io_sumIn_bits_last = PECross_124_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_125_multiply_io_input_io_sumOut_ready = PECross_126_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_125_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_125_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_125_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_125_multiply_io_input_io_actIn_valid = PECross_124_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_125_multiply_io_input_io_actIn_bits_x_0 = PECross_124_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_125_multiply_io_input_io_actIn_bits_last = PECross_124_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_125_multiply_io_input_io_weiIn_valid = PECross_109_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_125_multiply_io_input_io_weiIn_bits_x_0 = PECross_109_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_125_multiply_io_input_io_weiIn_bits_last = PECross_109_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_125_multiply_io_input_io_actOut_ready = PECross_126_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_125_multiply_io_input_io_weiOut_ready = PECross_141_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_126_clock = clock;
  assign PECross_126_reset = rst;
  assign PECross_126_multiply_io_input_io_sumIn_valid = PECross_125_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_126_multiply_io_input_io_sumIn_bits_x_0 = PECross_125_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_126_multiply_io_input_io_sumIn_bits_last = PECross_125_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_126_multiply_io_input_io_sumOut_ready = PECross_127_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_126_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_126_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_126_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_126_multiply_io_input_io_actIn_valid = PECross_125_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_126_multiply_io_input_io_actIn_bits_x_0 = PECross_125_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_126_multiply_io_input_io_actIn_bits_last = PECross_125_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_126_multiply_io_input_io_weiIn_valid = PECross_110_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_126_multiply_io_input_io_weiIn_bits_x_0 = PECross_110_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_126_multiply_io_input_io_weiIn_bits_last = PECross_110_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_126_multiply_io_input_io_actOut_ready = PECross_127_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_126_multiply_io_input_io_weiOut_ready = PECross_142_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_127_clock = clock;
  assign PECross_127_reset = rst;
  assign PECross_127_multiply_io_input_io_sumIn_valid = PECross_126_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_127_multiply_io_input_io_sumIn_bits_x_0 = PECross_126_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_127_multiply_io_input_io_sumIn_bits_last = PECross_126_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_127_multiply_io_input_io_sumOut_ready = io_sumOut_7_ready; // @[mac.scala 45:29]
  assign PECross_127_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_127_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_127_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_127_multiply_io_input_io_actIn_valid = PECross_126_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_127_multiply_io_input_io_actIn_bits_x_0 = PECross_126_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_127_multiply_io_input_io_actIn_bits_last = PECross_126_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_127_multiply_io_input_io_weiIn_valid = PECross_111_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_127_multiply_io_input_io_weiIn_bits_x_0 = PECross_111_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_127_multiply_io_input_io_weiIn_bits_last = PECross_111_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_127_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_127_multiply_io_input_io_weiOut_ready = PECross_143_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_128_clock = clock;
  assign PECross_128_reset = rst;
  assign PECross_128_multiply_io_input_io_sumIn_valid = io_sumIn_8_valid; // @[mac.scala 33:28]
  assign PECross_128_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_8_bits_x_0; // @[mac.scala 33:28]
  assign PECross_128_multiply_io_input_io_sumIn_bits_last = io_sumIn_8_bits_last; // @[mac.scala 33:28]
  assign PECross_128_multiply_io_input_io_sumOut_ready = PECross_129_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_128_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_128_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_128_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_128_multiply_io_input_io_actIn_valid = io_actIn_8_valid; // @[mac.scala 32:28]
  assign PECross_128_multiply_io_input_io_actIn_bits_x_0 = io_actIn_8_bits_x_0; // @[mac.scala 32:28]
  assign PECross_128_multiply_io_input_io_actIn_bits_last = io_actIn_8_bits_last; // @[mac.scala 32:28]
  assign PECross_128_multiply_io_input_io_weiIn_valid = PECross_112_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_128_multiply_io_input_io_weiIn_bits_x_0 = PECross_112_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_128_multiply_io_input_io_weiIn_bits_last = PECross_112_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_128_multiply_io_input_io_actOut_ready = PECross_129_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_128_multiply_io_input_io_weiOut_ready = PECross_144_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_129_clock = clock;
  assign PECross_129_reset = rst;
  assign PECross_129_multiply_io_input_io_sumIn_valid = PECross_128_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_129_multiply_io_input_io_sumIn_bits_x_0 = PECross_128_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_129_multiply_io_input_io_sumIn_bits_last = PECross_128_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_129_multiply_io_input_io_sumOut_ready = PECross_130_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_129_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_129_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_129_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_129_multiply_io_input_io_actIn_valid = PECross_128_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_129_multiply_io_input_io_actIn_bits_x_0 = PECross_128_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_129_multiply_io_input_io_actIn_bits_last = PECross_128_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_129_multiply_io_input_io_weiIn_valid = PECross_113_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_129_multiply_io_input_io_weiIn_bits_x_0 = PECross_113_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_129_multiply_io_input_io_weiIn_bits_last = PECross_113_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_129_multiply_io_input_io_actOut_ready = PECross_130_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_129_multiply_io_input_io_weiOut_ready = PECross_145_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_130_clock = clock;
  assign PECross_130_reset = rst;
  assign PECross_130_multiply_io_input_io_sumIn_valid = PECross_129_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_130_multiply_io_input_io_sumIn_bits_x_0 = PECross_129_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_130_multiply_io_input_io_sumIn_bits_last = PECross_129_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_130_multiply_io_input_io_sumOut_ready = PECross_131_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_130_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_130_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_130_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_130_multiply_io_input_io_actIn_valid = PECross_129_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_130_multiply_io_input_io_actIn_bits_x_0 = PECross_129_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_130_multiply_io_input_io_actIn_bits_last = PECross_129_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_130_multiply_io_input_io_weiIn_valid = PECross_114_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_130_multiply_io_input_io_weiIn_bits_x_0 = PECross_114_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_130_multiply_io_input_io_weiIn_bits_last = PECross_114_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_130_multiply_io_input_io_actOut_ready = PECross_131_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_130_multiply_io_input_io_weiOut_ready = PECross_146_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_131_clock = clock;
  assign PECross_131_reset = rst;
  assign PECross_131_multiply_io_input_io_sumIn_valid = PECross_130_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_131_multiply_io_input_io_sumIn_bits_x_0 = PECross_130_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_131_multiply_io_input_io_sumIn_bits_last = PECross_130_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_131_multiply_io_input_io_sumOut_ready = PECross_132_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_131_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_131_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_131_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_131_multiply_io_input_io_actIn_valid = PECross_130_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_131_multiply_io_input_io_actIn_bits_x_0 = PECross_130_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_131_multiply_io_input_io_actIn_bits_last = PECross_130_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_131_multiply_io_input_io_weiIn_valid = PECross_115_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_131_multiply_io_input_io_weiIn_bits_x_0 = PECross_115_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_131_multiply_io_input_io_weiIn_bits_last = PECross_115_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_131_multiply_io_input_io_actOut_ready = PECross_132_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_131_multiply_io_input_io_weiOut_ready = PECross_147_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_132_clock = clock;
  assign PECross_132_reset = rst;
  assign PECross_132_multiply_io_input_io_sumIn_valid = PECross_131_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_132_multiply_io_input_io_sumIn_bits_x_0 = PECross_131_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_132_multiply_io_input_io_sumIn_bits_last = PECross_131_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_132_multiply_io_input_io_sumOut_ready = PECross_133_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_132_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_132_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_132_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_132_multiply_io_input_io_actIn_valid = PECross_131_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_132_multiply_io_input_io_actIn_bits_x_0 = PECross_131_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_132_multiply_io_input_io_actIn_bits_last = PECross_131_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_132_multiply_io_input_io_weiIn_valid = PECross_116_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_132_multiply_io_input_io_weiIn_bits_x_0 = PECross_116_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_132_multiply_io_input_io_weiIn_bits_last = PECross_116_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_132_multiply_io_input_io_actOut_ready = PECross_133_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_132_multiply_io_input_io_weiOut_ready = PECross_148_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_133_clock = clock;
  assign PECross_133_reset = rst;
  assign PECross_133_multiply_io_input_io_sumIn_valid = PECross_132_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_133_multiply_io_input_io_sumIn_bits_x_0 = PECross_132_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_133_multiply_io_input_io_sumIn_bits_last = PECross_132_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_133_multiply_io_input_io_sumOut_ready = PECross_134_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_133_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_133_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_133_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_133_multiply_io_input_io_actIn_valid = PECross_132_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_133_multiply_io_input_io_actIn_bits_x_0 = PECross_132_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_133_multiply_io_input_io_actIn_bits_last = PECross_132_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_133_multiply_io_input_io_weiIn_valid = PECross_117_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_133_multiply_io_input_io_weiIn_bits_x_0 = PECross_117_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_133_multiply_io_input_io_weiIn_bits_last = PECross_117_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_133_multiply_io_input_io_actOut_ready = PECross_134_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_133_multiply_io_input_io_weiOut_ready = PECross_149_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_134_clock = clock;
  assign PECross_134_reset = rst;
  assign PECross_134_multiply_io_input_io_sumIn_valid = PECross_133_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_134_multiply_io_input_io_sumIn_bits_x_0 = PECross_133_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_134_multiply_io_input_io_sumIn_bits_last = PECross_133_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_134_multiply_io_input_io_sumOut_ready = PECross_135_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_134_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_134_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_134_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_134_multiply_io_input_io_actIn_valid = PECross_133_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_134_multiply_io_input_io_actIn_bits_x_0 = PECross_133_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_134_multiply_io_input_io_actIn_bits_last = PECross_133_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_134_multiply_io_input_io_weiIn_valid = PECross_118_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_134_multiply_io_input_io_weiIn_bits_x_0 = PECross_118_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_134_multiply_io_input_io_weiIn_bits_last = PECross_118_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_134_multiply_io_input_io_actOut_ready = PECross_135_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_134_multiply_io_input_io_weiOut_ready = PECross_150_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_135_clock = clock;
  assign PECross_135_reset = rst;
  assign PECross_135_multiply_io_input_io_sumIn_valid = PECross_134_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_135_multiply_io_input_io_sumIn_bits_x_0 = PECross_134_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_135_multiply_io_input_io_sumIn_bits_last = PECross_134_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_135_multiply_io_input_io_sumOut_ready = PECross_136_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_135_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_135_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_135_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_135_multiply_io_input_io_actIn_valid = PECross_134_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_135_multiply_io_input_io_actIn_bits_x_0 = PECross_134_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_135_multiply_io_input_io_actIn_bits_last = PECross_134_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_135_multiply_io_input_io_weiIn_valid = PECross_119_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_135_multiply_io_input_io_weiIn_bits_x_0 = PECross_119_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_135_multiply_io_input_io_weiIn_bits_last = PECross_119_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_135_multiply_io_input_io_actOut_ready = PECross_136_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_135_multiply_io_input_io_weiOut_ready = PECross_151_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_136_clock = clock;
  assign PECross_136_reset = rst;
  assign PECross_136_multiply_io_input_io_sumIn_valid = PECross_135_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_136_multiply_io_input_io_sumIn_bits_x_0 = PECross_135_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_136_multiply_io_input_io_sumIn_bits_last = PECross_135_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_136_multiply_io_input_io_sumOut_ready = PECross_137_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_136_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_136_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_136_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_136_multiply_io_input_io_actIn_valid = PECross_135_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_136_multiply_io_input_io_actIn_bits_x_0 = PECross_135_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_136_multiply_io_input_io_actIn_bits_last = PECross_135_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_136_multiply_io_input_io_weiIn_valid = PECross_120_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_136_multiply_io_input_io_weiIn_bits_x_0 = PECross_120_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_136_multiply_io_input_io_weiIn_bits_last = PECross_120_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_136_multiply_io_input_io_actOut_ready = PECross_137_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_136_multiply_io_input_io_weiOut_ready = PECross_152_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_137_clock = clock;
  assign PECross_137_reset = rst;
  assign PECross_137_multiply_io_input_io_sumIn_valid = PECross_136_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_137_multiply_io_input_io_sumIn_bits_x_0 = PECross_136_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_137_multiply_io_input_io_sumIn_bits_last = PECross_136_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_137_multiply_io_input_io_sumOut_ready = PECross_138_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_137_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_137_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_137_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_137_multiply_io_input_io_actIn_valid = PECross_136_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_137_multiply_io_input_io_actIn_bits_x_0 = PECross_136_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_137_multiply_io_input_io_actIn_bits_last = PECross_136_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_137_multiply_io_input_io_weiIn_valid = PECross_121_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_137_multiply_io_input_io_weiIn_bits_x_0 = PECross_121_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_137_multiply_io_input_io_weiIn_bits_last = PECross_121_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_137_multiply_io_input_io_actOut_ready = PECross_138_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_137_multiply_io_input_io_weiOut_ready = PECross_153_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_138_clock = clock;
  assign PECross_138_reset = rst;
  assign PECross_138_multiply_io_input_io_sumIn_valid = PECross_137_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_138_multiply_io_input_io_sumIn_bits_x_0 = PECross_137_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_138_multiply_io_input_io_sumIn_bits_last = PECross_137_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_138_multiply_io_input_io_sumOut_ready = PECross_139_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_138_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_138_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_138_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_138_multiply_io_input_io_actIn_valid = PECross_137_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_138_multiply_io_input_io_actIn_bits_x_0 = PECross_137_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_138_multiply_io_input_io_actIn_bits_last = PECross_137_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_138_multiply_io_input_io_weiIn_valid = PECross_122_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_138_multiply_io_input_io_weiIn_bits_x_0 = PECross_122_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_138_multiply_io_input_io_weiIn_bits_last = PECross_122_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_138_multiply_io_input_io_actOut_ready = PECross_139_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_138_multiply_io_input_io_weiOut_ready = PECross_154_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_139_clock = clock;
  assign PECross_139_reset = rst;
  assign PECross_139_multiply_io_input_io_sumIn_valid = PECross_138_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_139_multiply_io_input_io_sumIn_bits_x_0 = PECross_138_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_139_multiply_io_input_io_sumIn_bits_last = PECross_138_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_139_multiply_io_input_io_sumOut_ready = PECross_140_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_139_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_139_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_139_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_139_multiply_io_input_io_actIn_valid = PECross_138_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_139_multiply_io_input_io_actIn_bits_x_0 = PECross_138_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_139_multiply_io_input_io_actIn_bits_last = PECross_138_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_139_multiply_io_input_io_weiIn_valid = PECross_123_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_139_multiply_io_input_io_weiIn_bits_x_0 = PECross_123_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_139_multiply_io_input_io_weiIn_bits_last = PECross_123_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_139_multiply_io_input_io_actOut_ready = PECross_140_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_139_multiply_io_input_io_weiOut_ready = PECross_155_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_140_clock = clock;
  assign PECross_140_reset = rst;
  assign PECross_140_multiply_io_input_io_sumIn_valid = PECross_139_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_140_multiply_io_input_io_sumIn_bits_x_0 = PECross_139_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_140_multiply_io_input_io_sumIn_bits_last = PECross_139_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_140_multiply_io_input_io_sumOut_ready = PECross_141_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_140_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_140_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_140_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_140_multiply_io_input_io_actIn_valid = PECross_139_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_140_multiply_io_input_io_actIn_bits_x_0 = PECross_139_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_140_multiply_io_input_io_actIn_bits_last = PECross_139_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_140_multiply_io_input_io_weiIn_valid = PECross_124_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_140_multiply_io_input_io_weiIn_bits_x_0 = PECross_124_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_140_multiply_io_input_io_weiIn_bits_last = PECross_124_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_140_multiply_io_input_io_actOut_ready = PECross_141_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_140_multiply_io_input_io_weiOut_ready = PECross_156_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_141_clock = clock;
  assign PECross_141_reset = rst;
  assign PECross_141_multiply_io_input_io_sumIn_valid = PECross_140_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_141_multiply_io_input_io_sumIn_bits_x_0 = PECross_140_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_141_multiply_io_input_io_sumIn_bits_last = PECross_140_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_141_multiply_io_input_io_sumOut_ready = PECross_142_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_141_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_141_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_141_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_141_multiply_io_input_io_actIn_valid = PECross_140_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_141_multiply_io_input_io_actIn_bits_x_0 = PECross_140_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_141_multiply_io_input_io_actIn_bits_last = PECross_140_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_141_multiply_io_input_io_weiIn_valid = PECross_125_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_141_multiply_io_input_io_weiIn_bits_x_0 = PECross_125_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_141_multiply_io_input_io_weiIn_bits_last = PECross_125_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_141_multiply_io_input_io_actOut_ready = PECross_142_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_141_multiply_io_input_io_weiOut_ready = PECross_157_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_142_clock = clock;
  assign PECross_142_reset = rst;
  assign PECross_142_multiply_io_input_io_sumIn_valid = PECross_141_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_142_multiply_io_input_io_sumIn_bits_x_0 = PECross_141_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_142_multiply_io_input_io_sumIn_bits_last = PECross_141_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_142_multiply_io_input_io_sumOut_ready = PECross_143_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_142_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_142_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_142_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_142_multiply_io_input_io_actIn_valid = PECross_141_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_142_multiply_io_input_io_actIn_bits_x_0 = PECross_141_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_142_multiply_io_input_io_actIn_bits_last = PECross_141_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_142_multiply_io_input_io_weiIn_valid = PECross_126_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_142_multiply_io_input_io_weiIn_bits_x_0 = PECross_126_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_142_multiply_io_input_io_weiIn_bits_last = PECross_126_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_142_multiply_io_input_io_actOut_ready = PECross_143_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_142_multiply_io_input_io_weiOut_ready = PECross_158_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_143_clock = clock;
  assign PECross_143_reset = rst;
  assign PECross_143_multiply_io_input_io_sumIn_valid = PECross_142_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_143_multiply_io_input_io_sumIn_bits_x_0 = PECross_142_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_143_multiply_io_input_io_sumIn_bits_last = PECross_142_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_143_multiply_io_input_io_sumOut_ready = io_sumOut_8_ready; // @[mac.scala 45:29]
  assign PECross_143_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_143_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_143_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_143_multiply_io_input_io_actIn_valid = PECross_142_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_143_multiply_io_input_io_actIn_bits_x_0 = PECross_142_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_143_multiply_io_input_io_actIn_bits_last = PECross_142_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_143_multiply_io_input_io_weiIn_valid = PECross_127_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_143_multiply_io_input_io_weiIn_bits_x_0 = PECross_127_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_143_multiply_io_input_io_weiIn_bits_last = PECross_127_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_143_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_143_multiply_io_input_io_weiOut_ready = PECross_159_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_144_clock = clock;
  assign PECross_144_reset = rst;
  assign PECross_144_multiply_io_input_io_sumIn_valid = io_sumIn_9_valid; // @[mac.scala 33:28]
  assign PECross_144_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_9_bits_x_0; // @[mac.scala 33:28]
  assign PECross_144_multiply_io_input_io_sumIn_bits_last = io_sumIn_9_bits_last; // @[mac.scala 33:28]
  assign PECross_144_multiply_io_input_io_sumOut_ready = PECross_145_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_144_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_144_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_144_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_144_multiply_io_input_io_actIn_valid = io_actIn_9_valid; // @[mac.scala 32:28]
  assign PECross_144_multiply_io_input_io_actIn_bits_x_0 = io_actIn_9_bits_x_0; // @[mac.scala 32:28]
  assign PECross_144_multiply_io_input_io_actIn_bits_last = io_actIn_9_bits_last; // @[mac.scala 32:28]
  assign PECross_144_multiply_io_input_io_weiIn_valid = PECross_128_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_144_multiply_io_input_io_weiIn_bits_x_0 = PECross_128_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_144_multiply_io_input_io_weiIn_bits_last = PECross_128_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_144_multiply_io_input_io_actOut_ready = PECross_145_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_144_multiply_io_input_io_weiOut_ready = PECross_160_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_145_clock = clock;
  assign PECross_145_reset = rst;
  assign PECross_145_multiply_io_input_io_sumIn_valid = PECross_144_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_145_multiply_io_input_io_sumIn_bits_x_0 = PECross_144_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_145_multiply_io_input_io_sumIn_bits_last = PECross_144_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_145_multiply_io_input_io_sumOut_ready = PECross_146_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_145_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_145_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_145_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_145_multiply_io_input_io_actIn_valid = PECross_144_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_145_multiply_io_input_io_actIn_bits_x_0 = PECross_144_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_145_multiply_io_input_io_actIn_bits_last = PECross_144_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_145_multiply_io_input_io_weiIn_valid = PECross_129_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_145_multiply_io_input_io_weiIn_bits_x_0 = PECross_129_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_145_multiply_io_input_io_weiIn_bits_last = PECross_129_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_145_multiply_io_input_io_actOut_ready = PECross_146_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_145_multiply_io_input_io_weiOut_ready = PECross_161_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_146_clock = clock;
  assign PECross_146_reset = rst;
  assign PECross_146_multiply_io_input_io_sumIn_valid = PECross_145_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_146_multiply_io_input_io_sumIn_bits_x_0 = PECross_145_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_146_multiply_io_input_io_sumIn_bits_last = PECross_145_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_146_multiply_io_input_io_sumOut_ready = PECross_147_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_146_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_146_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_146_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_146_multiply_io_input_io_actIn_valid = PECross_145_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_146_multiply_io_input_io_actIn_bits_x_0 = PECross_145_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_146_multiply_io_input_io_actIn_bits_last = PECross_145_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_146_multiply_io_input_io_weiIn_valid = PECross_130_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_146_multiply_io_input_io_weiIn_bits_x_0 = PECross_130_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_146_multiply_io_input_io_weiIn_bits_last = PECross_130_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_146_multiply_io_input_io_actOut_ready = PECross_147_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_146_multiply_io_input_io_weiOut_ready = PECross_162_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_147_clock = clock;
  assign PECross_147_reset = rst;
  assign PECross_147_multiply_io_input_io_sumIn_valid = PECross_146_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_147_multiply_io_input_io_sumIn_bits_x_0 = PECross_146_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_147_multiply_io_input_io_sumIn_bits_last = PECross_146_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_147_multiply_io_input_io_sumOut_ready = PECross_148_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_147_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_147_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_147_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_147_multiply_io_input_io_actIn_valid = PECross_146_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_147_multiply_io_input_io_actIn_bits_x_0 = PECross_146_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_147_multiply_io_input_io_actIn_bits_last = PECross_146_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_147_multiply_io_input_io_weiIn_valid = PECross_131_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_147_multiply_io_input_io_weiIn_bits_x_0 = PECross_131_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_147_multiply_io_input_io_weiIn_bits_last = PECross_131_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_147_multiply_io_input_io_actOut_ready = PECross_148_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_147_multiply_io_input_io_weiOut_ready = PECross_163_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_148_clock = clock;
  assign PECross_148_reset = rst;
  assign PECross_148_multiply_io_input_io_sumIn_valid = PECross_147_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_148_multiply_io_input_io_sumIn_bits_x_0 = PECross_147_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_148_multiply_io_input_io_sumIn_bits_last = PECross_147_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_148_multiply_io_input_io_sumOut_ready = PECross_149_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_148_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_148_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_148_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_148_multiply_io_input_io_actIn_valid = PECross_147_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_148_multiply_io_input_io_actIn_bits_x_0 = PECross_147_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_148_multiply_io_input_io_actIn_bits_last = PECross_147_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_148_multiply_io_input_io_weiIn_valid = PECross_132_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_148_multiply_io_input_io_weiIn_bits_x_0 = PECross_132_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_148_multiply_io_input_io_weiIn_bits_last = PECross_132_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_148_multiply_io_input_io_actOut_ready = PECross_149_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_148_multiply_io_input_io_weiOut_ready = PECross_164_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_149_clock = clock;
  assign PECross_149_reset = rst;
  assign PECross_149_multiply_io_input_io_sumIn_valid = PECross_148_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_149_multiply_io_input_io_sumIn_bits_x_0 = PECross_148_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_149_multiply_io_input_io_sumIn_bits_last = PECross_148_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_149_multiply_io_input_io_sumOut_ready = PECross_150_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_149_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_149_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_149_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_149_multiply_io_input_io_actIn_valid = PECross_148_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_149_multiply_io_input_io_actIn_bits_x_0 = PECross_148_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_149_multiply_io_input_io_actIn_bits_last = PECross_148_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_149_multiply_io_input_io_weiIn_valid = PECross_133_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_149_multiply_io_input_io_weiIn_bits_x_0 = PECross_133_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_149_multiply_io_input_io_weiIn_bits_last = PECross_133_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_149_multiply_io_input_io_actOut_ready = PECross_150_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_149_multiply_io_input_io_weiOut_ready = PECross_165_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_150_clock = clock;
  assign PECross_150_reset = rst;
  assign PECross_150_multiply_io_input_io_sumIn_valid = PECross_149_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_150_multiply_io_input_io_sumIn_bits_x_0 = PECross_149_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_150_multiply_io_input_io_sumIn_bits_last = PECross_149_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_150_multiply_io_input_io_sumOut_ready = PECross_151_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_150_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_150_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_150_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_150_multiply_io_input_io_actIn_valid = PECross_149_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_150_multiply_io_input_io_actIn_bits_x_0 = PECross_149_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_150_multiply_io_input_io_actIn_bits_last = PECross_149_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_150_multiply_io_input_io_weiIn_valid = PECross_134_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_150_multiply_io_input_io_weiIn_bits_x_0 = PECross_134_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_150_multiply_io_input_io_weiIn_bits_last = PECross_134_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_150_multiply_io_input_io_actOut_ready = PECross_151_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_150_multiply_io_input_io_weiOut_ready = PECross_166_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_151_clock = clock;
  assign PECross_151_reset = rst;
  assign PECross_151_multiply_io_input_io_sumIn_valid = PECross_150_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_151_multiply_io_input_io_sumIn_bits_x_0 = PECross_150_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_151_multiply_io_input_io_sumIn_bits_last = PECross_150_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_151_multiply_io_input_io_sumOut_ready = PECross_152_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_151_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_151_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_151_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_151_multiply_io_input_io_actIn_valid = PECross_150_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_151_multiply_io_input_io_actIn_bits_x_0 = PECross_150_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_151_multiply_io_input_io_actIn_bits_last = PECross_150_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_151_multiply_io_input_io_weiIn_valid = PECross_135_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_151_multiply_io_input_io_weiIn_bits_x_0 = PECross_135_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_151_multiply_io_input_io_weiIn_bits_last = PECross_135_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_151_multiply_io_input_io_actOut_ready = PECross_152_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_151_multiply_io_input_io_weiOut_ready = PECross_167_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_152_clock = clock;
  assign PECross_152_reset = rst;
  assign PECross_152_multiply_io_input_io_sumIn_valid = PECross_151_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_152_multiply_io_input_io_sumIn_bits_x_0 = PECross_151_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_152_multiply_io_input_io_sumIn_bits_last = PECross_151_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_152_multiply_io_input_io_sumOut_ready = PECross_153_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_152_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_152_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_152_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_152_multiply_io_input_io_actIn_valid = PECross_151_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_152_multiply_io_input_io_actIn_bits_x_0 = PECross_151_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_152_multiply_io_input_io_actIn_bits_last = PECross_151_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_152_multiply_io_input_io_weiIn_valid = PECross_136_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_152_multiply_io_input_io_weiIn_bits_x_0 = PECross_136_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_152_multiply_io_input_io_weiIn_bits_last = PECross_136_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_152_multiply_io_input_io_actOut_ready = PECross_153_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_152_multiply_io_input_io_weiOut_ready = PECross_168_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_153_clock = clock;
  assign PECross_153_reset = rst;
  assign PECross_153_multiply_io_input_io_sumIn_valid = PECross_152_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_153_multiply_io_input_io_sumIn_bits_x_0 = PECross_152_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_153_multiply_io_input_io_sumIn_bits_last = PECross_152_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_153_multiply_io_input_io_sumOut_ready = PECross_154_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_153_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_153_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_153_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_153_multiply_io_input_io_actIn_valid = PECross_152_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_153_multiply_io_input_io_actIn_bits_x_0 = PECross_152_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_153_multiply_io_input_io_actIn_bits_last = PECross_152_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_153_multiply_io_input_io_weiIn_valid = PECross_137_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_153_multiply_io_input_io_weiIn_bits_x_0 = PECross_137_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_153_multiply_io_input_io_weiIn_bits_last = PECross_137_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_153_multiply_io_input_io_actOut_ready = PECross_154_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_153_multiply_io_input_io_weiOut_ready = PECross_169_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_154_clock = clock;
  assign PECross_154_reset = rst;
  assign PECross_154_multiply_io_input_io_sumIn_valid = PECross_153_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_154_multiply_io_input_io_sumIn_bits_x_0 = PECross_153_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_154_multiply_io_input_io_sumIn_bits_last = PECross_153_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_154_multiply_io_input_io_sumOut_ready = PECross_155_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_154_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_154_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_154_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_154_multiply_io_input_io_actIn_valid = PECross_153_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_154_multiply_io_input_io_actIn_bits_x_0 = PECross_153_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_154_multiply_io_input_io_actIn_bits_last = PECross_153_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_154_multiply_io_input_io_weiIn_valid = PECross_138_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_154_multiply_io_input_io_weiIn_bits_x_0 = PECross_138_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_154_multiply_io_input_io_weiIn_bits_last = PECross_138_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_154_multiply_io_input_io_actOut_ready = PECross_155_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_154_multiply_io_input_io_weiOut_ready = PECross_170_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_155_clock = clock;
  assign PECross_155_reset = rst;
  assign PECross_155_multiply_io_input_io_sumIn_valid = PECross_154_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_155_multiply_io_input_io_sumIn_bits_x_0 = PECross_154_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_155_multiply_io_input_io_sumIn_bits_last = PECross_154_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_155_multiply_io_input_io_sumOut_ready = PECross_156_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_155_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_155_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_155_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_155_multiply_io_input_io_actIn_valid = PECross_154_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_155_multiply_io_input_io_actIn_bits_x_0 = PECross_154_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_155_multiply_io_input_io_actIn_bits_last = PECross_154_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_155_multiply_io_input_io_weiIn_valid = PECross_139_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_155_multiply_io_input_io_weiIn_bits_x_0 = PECross_139_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_155_multiply_io_input_io_weiIn_bits_last = PECross_139_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_155_multiply_io_input_io_actOut_ready = PECross_156_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_155_multiply_io_input_io_weiOut_ready = PECross_171_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_156_clock = clock;
  assign PECross_156_reset = rst;
  assign PECross_156_multiply_io_input_io_sumIn_valid = PECross_155_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_156_multiply_io_input_io_sumIn_bits_x_0 = PECross_155_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_156_multiply_io_input_io_sumIn_bits_last = PECross_155_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_156_multiply_io_input_io_sumOut_ready = PECross_157_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_156_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_156_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_156_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_156_multiply_io_input_io_actIn_valid = PECross_155_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_156_multiply_io_input_io_actIn_bits_x_0 = PECross_155_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_156_multiply_io_input_io_actIn_bits_last = PECross_155_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_156_multiply_io_input_io_weiIn_valid = PECross_140_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_156_multiply_io_input_io_weiIn_bits_x_0 = PECross_140_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_156_multiply_io_input_io_weiIn_bits_last = PECross_140_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_156_multiply_io_input_io_actOut_ready = PECross_157_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_156_multiply_io_input_io_weiOut_ready = PECross_172_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_157_clock = clock;
  assign PECross_157_reset = rst;
  assign PECross_157_multiply_io_input_io_sumIn_valid = PECross_156_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_157_multiply_io_input_io_sumIn_bits_x_0 = PECross_156_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_157_multiply_io_input_io_sumIn_bits_last = PECross_156_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_157_multiply_io_input_io_sumOut_ready = PECross_158_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_157_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_157_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_157_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_157_multiply_io_input_io_actIn_valid = PECross_156_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_157_multiply_io_input_io_actIn_bits_x_0 = PECross_156_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_157_multiply_io_input_io_actIn_bits_last = PECross_156_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_157_multiply_io_input_io_weiIn_valid = PECross_141_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_157_multiply_io_input_io_weiIn_bits_x_0 = PECross_141_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_157_multiply_io_input_io_weiIn_bits_last = PECross_141_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_157_multiply_io_input_io_actOut_ready = PECross_158_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_157_multiply_io_input_io_weiOut_ready = PECross_173_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_158_clock = clock;
  assign PECross_158_reset = rst;
  assign PECross_158_multiply_io_input_io_sumIn_valid = PECross_157_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_158_multiply_io_input_io_sumIn_bits_x_0 = PECross_157_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_158_multiply_io_input_io_sumIn_bits_last = PECross_157_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_158_multiply_io_input_io_sumOut_ready = PECross_159_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_158_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_158_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_158_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_158_multiply_io_input_io_actIn_valid = PECross_157_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_158_multiply_io_input_io_actIn_bits_x_0 = PECross_157_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_158_multiply_io_input_io_actIn_bits_last = PECross_157_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_158_multiply_io_input_io_weiIn_valid = PECross_142_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_158_multiply_io_input_io_weiIn_bits_x_0 = PECross_142_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_158_multiply_io_input_io_weiIn_bits_last = PECross_142_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_158_multiply_io_input_io_actOut_ready = PECross_159_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_158_multiply_io_input_io_weiOut_ready = PECross_174_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_159_clock = clock;
  assign PECross_159_reset = rst;
  assign PECross_159_multiply_io_input_io_sumIn_valid = PECross_158_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_159_multiply_io_input_io_sumIn_bits_x_0 = PECross_158_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_159_multiply_io_input_io_sumIn_bits_last = PECross_158_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_159_multiply_io_input_io_sumOut_ready = io_sumOut_9_ready; // @[mac.scala 45:29]
  assign PECross_159_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_159_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_159_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_159_multiply_io_input_io_actIn_valid = PECross_158_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_159_multiply_io_input_io_actIn_bits_x_0 = PECross_158_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_159_multiply_io_input_io_actIn_bits_last = PECross_158_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_159_multiply_io_input_io_weiIn_valid = PECross_143_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_159_multiply_io_input_io_weiIn_bits_x_0 = PECross_143_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_159_multiply_io_input_io_weiIn_bits_last = PECross_143_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_159_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_159_multiply_io_input_io_weiOut_ready = PECross_175_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_160_clock = clock;
  assign PECross_160_reset = rst;
  assign PECross_160_multiply_io_input_io_sumIn_valid = io_sumIn_10_valid; // @[mac.scala 33:28]
  assign PECross_160_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_10_bits_x_0; // @[mac.scala 33:28]
  assign PECross_160_multiply_io_input_io_sumIn_bits_last = io_sumIn_10_bits_last; // @[mac.scala 33:28]
  assign PECross_160_multiply_io_input_io_sumOut_ready = PECross_161_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_160_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_160_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_160_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_160_multiply_io_input_io_actIn_valid = io_actIn_10_valid; // @[mac.scala 32:28]
  assign PECross_160_multiply_io_input_io_actIn_bits_x_0 = io_actIn_10_bits_x_0; // @[mac.scala 32:28]
  assign PECross_160_multiply_io_input_io_actIn_bits_last = io_actIn_10_bits_last; // @[mac.scala 32:28]
  assign PECross_160_multiply_io_input_io_weiIn_valid = PECross_144_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_160_multiply_io_input_io_weiIn_bits_x_0 = PECross_144_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_160_multiply_io_input_io_weiIn_bits_last = PECross_144_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_160_multiply_io_input_io_actOut_ready = PECross_161_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_160_multiply_io_input_io_weiOut_ready = PECross_176_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_161_clock = clock;
  assign PECross_161_reset = rst;
  assign PECross_161_multiply_io_input_io_sumIn_valid = PECross_160_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_161_multiply_io_input_io_sumIn_bits_x_0 = PECross_160_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_161_multiply_io_input_io_sumIn_bits_last = PECross_160_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_161_multiply_io_input_io_sumOut_ready = PECross_162_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_161_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_161_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_161_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_161_multiply_io_input_io_actIn_valid = PECross_160_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_161_multiply_io_input_io_actIn_bits_x_0 = PECross_160_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_161_multiply_io_input_io_actIn_bits_last = PECross_160_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_161_multiply_io_input_io_weiIn_valid = PECross_145_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_161_multiply_io_input_io_weiIn_bits_x_0 = PECross_145_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_161_multiply_io_input_io_weiIn_bits_last = PECross_145_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_161_multiply_io_input_io_actOut_ready = PECross_162_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_161_multiply_io_input_io_weiOut_ready = PECross_177_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_162_clock = clock;
  assign PECross_162_reset = rst;
  assign PECross_162_multiply_io_input_io_sumIn_valid = PECross_161_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_162_multiply_io_input_io_sumIn_bits_x_0 = PECross_161_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_162_multiply_io_input_io_sumIn_bits_last = PECross_161_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_162_multiply_io_input_io_sumOut_ready = PECross_163_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_162_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_162_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_162_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_162_multiply_io_input_io_actIn_valid = PECross_161_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_162_multiply_io_input_io_actIn_bits_x_0 = PECross_161_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_162_multiply_io_input_io_actIn_bits_last = PECross_161_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_162_multiply_io_input_io_weiIn_valid = PECross_146_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_162_multiply_io_input_io_weiIn_bits_x_0 = PECross_146_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_162_multiply_io_input_io_weiIn_bits_last = PECross_146_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_162_multiply_io_input_io_actOut_ready = PECross_163_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_162_multiply_io_input_io_weiOut_ready = PECross_178_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_163_clock = clock;
  assign PECross_163_reset = rst;
  assign PECross_163_multiply_io_input_io_sumIn_valid = PECross_162_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_163_multiply_io_input_io_sumIn_bits_x_0 = PECross_162_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_163_multiply_io_input_io_sumIn_bits_last = PECross_162_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_163_multiply_io_input_io_sumOut_ready = PECross_164_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_163_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_163_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_163_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_163_multiply_io_input_io_actIn_valid = PECross_162_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_163_multiply_io_input_io_actIn_bits_x_0 = PECross_162_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_163_multiply_io_input_io_actIn_bits_last = PECross_162_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_163_multiply_io_input_io_weiIn_valid = PECross_147_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_163_multiply_io_input_io_weiIn_bits_x_0 = PECross_147_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_163_multiply_io_input_io_weiIn_bits_last = PECross_147_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_163_multiply_io_input_io_actOut_ready = PECross_164_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_163_multiply_io_input_io_weiOut_ready = PECross_179_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_164_clock = clock;
  assign PECross_164_reset = rst;
  assign PECross_164_multiply_io_input_io_sumIn_valid = PECross_163_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_164_multiply_io_input_io_sumIn_bits_x_0 = PECross_163_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_164_multiply_io_input_io_sumIn_bits_last = PECross_163_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_164_multiply_io_input_io_sumOut_ready = PECross_165_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_164_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_164_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_164_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_164_multiply_io_input_io_actIn_valid = PECross_163_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_164_multiply_io_input_io_actIn_bits_x_0 = PECross_163_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_164_multiply_io_input_io_actIn_bits_last = PECross_163_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_164_multiply_io_input_io_weiIn_valid = PECross_148_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_164_multiply_io_input_io_weiIn_bits_x_0 = PECross_148_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_164_multiply_io_input_io_weiIn_bits_last = PECross_148_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_164_multiply_io_input_io_actOut_ready = PECross_165_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_164_multiply_io_input_io_weiOut_ready = PECross_180_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_165_clock = clock;
  assign PECross_165_reset = rst;
  assign PECross_165_multiply_io_input_io_sumIn_valid = PECross_164_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_165_multiply_io_input_io_sumIn_bits_x_0 = PECross_164_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_165_multiply_io_input_io_sumIn_bits_last = PECross_164_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_165_multiply_io_input_io_sumOut_ready = PECross_166_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_165_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_165_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_165_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_165_multiply_io_input_io_actIn_valid = PECross_164_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_165_multiply_io_input_io_actIn_bits_x_0 = PECross_164_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_165_multiply_io_input_io_actIn_bits_last = PECross_164_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_165_multiply_io_input_io_weiIn_valid = PECross_149_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_165_multiply_io_input_io_weiIn_bits_x_0 = PECross_149_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_165_multiply_io_input_io_weiIn_bits_last = PECross_149_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_165_multiply_io_input_io_actOut_ready = PECross_166_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_165_multiply_io_input_io_weiOut_ready = PECross_181_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_166_clock = clock;
  assign PECross_166_reset = rst;
  assign PECross_166_multiply_io_input_io_sumIn_valid = PECross_165_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_166_multiply_io_input_io_sumIn_bits_x_0 = PECross_165_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_166_multiply_io_input_io_sumIn_bits_last = PECross_165_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_166_multiply_io_input_io_sumOut_ready = PECross_167_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_166_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_166_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_166_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_166_multiply_io_input_io_actIn_valid = PECross_165_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_166_multiply_io_input_io_actIn_bits_x_0 = PECross_165_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_166_multiply_io_input_io_actIn_bits_last = PECross_165_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_166_multiply_io_input_io_weiIn_valid = PECross_150_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_166_multiply_io_input_io_weiIn_bits_x_0 = PECross_150_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_166_multiply_io_input_io_weiIn_bits_last = PECross_150_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_166_multiply_io_input_io_actOut_ready = PECross_167_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_166_multiply_io_input_io_weiOut_ready = PECross_182_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_167_clock = clock;
  assign PECross_167_reset = rst;
  assign PECross_167_multiply_io_input_io_sumIn_valid = PECross_166_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_167_multiply_io_input_io_sumIn_bits_x_0 = PECross_166_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_167_multiply_io_input_io_sumIn_bits_last = PECross_166_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_167_multiply_io_input_io_sumOut_ready = PECross_168_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_167_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_167_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_167_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_167_multiply_io_input_io_actIn_valid = PECross_166_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_167_multiply_io_input_io_actIn_bits_x_0 = PECross_166_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_167_multiply_io_input_io_actIn_bits_last = PECross_166_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_167_multiply_io_input_io_weiIn_valid = PECross_151_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_167_multiply_io_input_io_weiIn_bits_x_0 = PECross_151_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_167_multiply_io_input_io_weiIn_bits_last = PECross_151_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_167_multiply_io_input_io_actOut_ready = PECross_168_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_167_multiply_io_input_io_weiOut_ready = PECross_183_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_168_clock = clock;
  assign PECross_168_reset = rst;
  assign PECross_168_multiply_io_input_io_sumIn_valid = PECross_167_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_168_multiply_io_input_io_sumIn_bits_x_0 = PECross_167_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_168_multiply_io_input_io_sumIn_bits_last = PECross_167_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_168_multiply_io_input_io_sumOut_ready = PECross_169_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_168_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_168_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_168_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_168_multiply_io_input_io_actIn_valid = PECross_167_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_168_multiply_io_input_io_actIn_bits_x_0 = PECross_167_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_168_multiply_io_input_io_actIn_bits_last = PECross_167_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_168_multiply_io_input_io_weiIn_valid = PECross_152_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_168_multiply_io_input_io_weiIn_bits_x_0 = PECross_152_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_168_multiply_io_input_io_weiIn_bits_last = PECross_152_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_168_multiply_io_input_io_actOut_ready = PECross_169_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_168_multiply_io_input_io_weiOut_ready = PECross_184_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_169_clock = clock;
  assign PECross_169_reset = rst;
  assign PECross_169_multiply_io_input_io_sumIn_valid = PECross_168_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_169_multiply_io_input_io_sumIn_bits_x_0 = PECross_168_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_169_multiply_io_input_io_sumIn_bits_last = PECross_168_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_169_multiply_io_input_io_sumOut_ready = PECross_170_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_169_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_169_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_169_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_169_multiply_io_input_io_actIn_valid = PECross_168_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_169_multiply_io_input_io_actIn_bits_x_0 = PECross_168_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_169_multiply_io_input_io_actIn_bits_last = PECross_168_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_169_multiply_io_input_io_weiIn_valid = PECross_153_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_169_multiply_io_input_io_weiIn_bits_x_0 = PECross_153_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_169_multiply_io_input_io_weiIn_bits_last = PECross_153_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_169_multiply_io_input_io_actOut_ready = PECross_170_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_169_multiply_io_input_io_weiOut_ready = PECross_185_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_170_clock = clock;
  assign PECross_170_reset = rst;
  assign PECross_170_multiply_io_input_io_sumIn_valid = PECross_169_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_170_multiply_io_input_io_sumIn_bits_x_0 = PECross_169_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_170_multiply_io_input_io_sumIn_bits_last = PECross_169_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_170_multiply_io_input_io_sumOut_ready = PECross_171_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_170_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_170_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_170_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_170_multiply_io_input_io_actIn_valid = PECross_169_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_170_multiply_io_input_io_actIn_bits_x_0 = PECross_169_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_170_multiply_io_input_io_actIn_bits_last = PECross_169_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_170_multiply_io_input_io_weiIn_valid = PECross_154_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_170_multiply_io_input_io_weiIn_bits_x_0 = PECross_154_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_170_multiply_io_input_io_weiIn_bits_last = PECross_154_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_170_multiply_io_input_io_actOut_ready = PECross_171_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_170_multiply_io_input_io_weiOut_ready = PECross_186_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_171_clock = clock;
  assign PECross_171_reset = rst;
  assign PECross_171_multiply_io_input_io_sumIn_valid = PECross_170_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_171_multiply_io_input_io_sumIn_bits_x_0 = PECross_170_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_171_multiply_io_input_io_sumIn_bits_last = PECross_170_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_171_multiply_io_input_io_sumOut_ready = PECross_172_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_171_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_171_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_171_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_171_multiply_io_input_io_actIn_valid = PECross_170_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_171_multiply_io_input_io_actIn_bits_x_0 = PECross_170_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_171_multiply_io_input_io_actIn_bits_last = PECross_170_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_171_multiply_io_input_io_weiIn_valid = PECross_155_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_171_multiply_io_input_io_weiIn_bits_x_0 = PECross_155_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_171_multiply_io_input_io_weiIn_bits_last = PECross_155_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_171_multiply_io_input_io_actOut_ready = PECross_172_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_171_multiply_io_input_io_weiOut_ready = PECross_187_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_172_clock = clock;
  assign PECross_172_reset = rst;
  assign PECross_172_multiply_io_input_io_sumIn_valid = PECross_171_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_172_multiply_io_input_io_sumIn_bits_x_0 = PECross_171_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_172_multiply_io_input_io_sumIn_bits_last = PECross_171_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_172_multiply_io_input_io_sumOut_ready = PECross_173_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_172_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_172_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_172_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_172_multiply_io_input_io_actIn_valid = PECross_171_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_172_multiply_io_input_io_actIn_bits_x_0 = PECross_171_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_172_multiply_io_input_io_actIn_bits_last = PECross_171_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_172_multiply_io_input_io_weiIn_valid = PECross_156_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_172_multiply_io_input_io_weiIn_bits_x_0 = PECross_156_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_172_multiply_io_input_io_weiIn_bits_last = PECross_156_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_172_multiply_io_input_io_actOut_ready = PECross_173_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_172_multiply_io_input_io_weiOut_ready = PECross_188_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_173_clock = clock;
  assign PECross_173_reset = rst;
  assign PECross_173_multiply_io_input_io_sumIn_valid = PECross_172_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_173_multiply_io_input_io_sumIn_bits_x_0 = PECross_172_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_173_multiply_io_input_io_sumIn_bits_last = PECross_172_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_173_multiply_io_input_io_sumOut_ready = PECross_174_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_173_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_173_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_173_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_173_multiply_io_input_io_actIn_valid = PECross_172_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_173_multiply_io_input_io_actIn_bits_x_0 = PECross_172_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_173_multiply_io_input_io_actIn_bits_last = PECross_172_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_173_multiply_io_input_io_weiIn_valid = PECross_157_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_173_multiply_io_input_io_weiIn_bits_x_0 = PECross_157_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_173_multiply_io_input_io_weiIn_bits_last = PECross_157_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_173_multiply_io_input_io_actOut_ready = PECross_174_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_173_multiply_io_input_io_weiOut_ready = PECross_189_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_174_clock = clock;
  assign PECross_174_reset = rst;
  assign PECross_174_multiply_io_input_io_sumIn_valid = PECross_173_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_174_multiply_io_input_io_sumIn_bits_x_0 = PECross_173_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_174_multiply_io_input_io_sumIn_bits_last = PECross_173_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_174_multiply_io_input_io_sumOut_ready = PECross_175_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_174_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_174_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_174_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_174_multiply_io_input_io_actIn_valid = PECross_173_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_174_multiply_io_input_io_actIn_bits_x_0 = PECross_173_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_174_multiply_io_input_io_actIn_bits_last = PECross_173_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_174_multiply_io_input_io_weiIn_valid = PECross_158_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_174_multiply_io_input_io_weiIn_bits_x_0 = PECross_158_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_174_multiply_io_input_io_weiIn_bits_last = PECross_158_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_174_multiply_io_input_io_actOut_ready = PECross_175_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_174_multiply_io_input_io_weiOut_ready = PECross_190_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_175_clock = clock;
  assign PECross_175_reset = rst;
  assign PECross_175_multiply_io_input_io_sumIn_valid = PECross_174_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_175_multiply_io_input_io_sumIn_bits_x_0 = PECross_174_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_175_multiply_io_input_io_sumIn_bits_last = PECross_174_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_175_multiply_io_input_io_sumOut_ready = io_sumOut_10_ready; // @[mac.scala 45:29]
  assign PECross_175_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_175_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_175_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_175_multiply_io_input_io_actIn_valid = PECross_174_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_175_multiply_io_input_io_actIn_bits_x_0 = PECross_174_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_175_multiply_io_input_io_actIn_bits_last = PECross_174_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_175_multiply_io_input_io_weiIn_valid = PECross_159_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_175_multiply_io_input_io_weiIn_bits_x_0 = PECross_159_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_175_multiply_io_input_io_weiIn_bits_last = PECross_159_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_175_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_175_multiply_io_input_io_weiOut_ready = PECross_191_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_176_clock = clock;
  assign PECross_176_reset = rst;
  assign PECross_176_multiply_io_input_io_sumIn_valid = io_sumIn_11_valid; // @[mac.scala 33:28]
  assign PECross_176_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_11_bits_x_0; // @[mac.scala 33:28]
  assign PECross_176_multiply_io_input_io_sumIn_bits_last = io_sumIn_11_bits_last; // @[mac.scala 33:28]
  assign PECross_176_multiply_io_input_io_sumOut_ready = PECross_177_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_176_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_176_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_176_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_176_multiply_io_input_io_actIn_valid = io_actIn_11_valid; // @[mac.scala 32:28]
  assign PECross_176_multiply_io_input_io_actIn_bits_x_0 = io_actIn_11_bits_x_0; // @[mac.scala 32:28]
  assign PECross_176_multiply_io_input_io_actIn_bits_last = io_actIn_11_bits_last; // @[mac.scala 32:28]
  assign PECross_176_multiply_io_input_io_weiIn_valid = PECross_160_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_176_multiply_io_input_io_weiIn_bits_x_0 = PECross_160_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_176_multiply_io_input_io_weiIn_bits_last = PECross_160_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_176_multiply_io_input_io_actOut_ready = PECross_177_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_176_multiply_io_input_io_weiOut_ready = PECross_192_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_177_clock = clock;
  assign PECross_177_reset = rst;
  assign PECross_177_multiply_io_input_io_sumIn_valid = PECross_176_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_177_multiply_io_input_io_sumIn_bits_x_0 = PECross_176_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_177_multiply_io_input_io_sumIn_bits_last = PECross_176_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_177_multiply_io_input_io_sumOut_ready = PECross_178_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_177_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_177_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_177_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_177_multiply_io_input_io_actIn_valid = PECross_176_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_177_multiply_io_input_io_actIn_bits_x_0 = PECross_176_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_177_multiply_io_input_io_actIn_bits_last = PECross_176_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_177_multiply_io_input_io_weiIn_valid = PECross_161_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_177_multiply_io_input_io_weiIn_bits_x_0 = PECross_161_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_177_multiply_io_input_io_weiIn_bits_last = PECross_161_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_177_multiply_io_input_io_actOut_ready = PECross_178_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_177_multiply_io_input_io_weiOut_ready = PECross_193_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_178_clock = clock;
  assign PECross_178_reset = rst;
  assign PECross_178_multiply_io_input_io_sumIn_valid = PECross_177_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_178_multiply_io_input_io_sumIn_bits_x_0 = PECross_177_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_178_multiply_io_input_io_sumIn_bits_last = PECross_177_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_178_multiply_io_input_io_sumOut_ready = PECross_179_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_178_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_178_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_178_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_178_multiply_io_input_io_actIn_valid = PECross_177_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_178_multiply_io_input_io_actIn_bits_x_0 = PECross_177_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_178_multiply_io_input_io_actIn_bits_last = PECross_177_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_178_multiply_io_input_io_weiIn_valid = PECross_162_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_178_multiply_io_input_io_weiIn_bits_x_0 = PECross_162_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_178_multiply_io_input_io_weiIn_bits_last = PECross_162_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_178_multiply_io_input_io_actOut_ready = PECross_179_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_178_multiply_io_input_io_weiOut_ready = PECross_194_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_179_clock = clock;
  assign PECross_179_reset = rst;
  assign PECross_179_multiply_io_input_io_sumIn_valid = PECross_178_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_179_multiply_io_input_io_sumIn_bits_x_0 = PECross_178_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_179_multiply_io_input_io_sumIn_bits_last = PECross_178_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_179_multiply_io_input_io_sumOut_ready = PECross_180_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_179_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_179_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_179_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_179_multiply_io_input_io_actIn_valid = PECross_178_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_179_multiply_io_input_io_actIn_bits_x_0 = PECross_178_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_179_multiply_io_input_io_actIn_bits_last = PECross_178_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_179_multiply_io_input_io_weiIn_valid = PECross_163_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_179_multiply_io_input_io_weiIn_bits_x_0 = PECross_163_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_179_multiply_io_input_io_weiIn_bits_last = PECross_163_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_179_multiply_io_input_io_actOut_ready = PECross_180_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_179_multiply_io_input_io_weiOut_ready = PECross_195_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_180_clock = clock;
  assign PECross_180_reset = rst;
  assign PECross_180_multiply_io_input_io_sumIn_valid = PECross_179_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_180_multiply_io_input_io_sumIn_bits_x_0 = PECross_179_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_180_multiply_io_input_io_sumIn_bits_last = PECross_179_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_180_multiply_io_input_io_sumOut_ready = PECross_181_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_180_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_180_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_180_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_180_multiply_io_input_io_actIn_valid = PECross_179_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_180_multiply_io_input_io_actIn_bits_x_0 = PECross_179_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_180_multiply_io_input_io_actIn_bits_last = PECross_179_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_180_multiply_io_input_io_weiIn_valid = PECross_164_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_180_multiply_io_input_io_weiIn_bits_x_0 = PECross_164_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_180_multiply_io_input_io_weiIn_bits_last = PECross_164_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_180_multiply_io_input_io_actOut_ready = PECross_181_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_180_multiply_io_input_io_weiOut_ready = PECross_196_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_181_clock = clock;
  assign PECross_181_reset = rst;
  assign PECross_181_multiply_io_input_io_sumIn_valid = PECross_180_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_181_multiply_io_input_io_sumIn_bits_x_0 = PECross_180_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_181_multiply_io_input_io_sumIn_bits_last = PECross_180_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_181_multiply_io_input_io_sumOut_ready = PECross_182_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_181_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_181_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_181_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_181_multiply_io_input_io_actIn_valid = PECross_180_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_181_multiply_io_input_io_actIn_bits_x_0 = PECross_180_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_181_multiply_io_input_io_actIn_bits_last = PECross_180_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_181_multiply_io_input_io_weiIn_valid = PECross_165_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_181_multiply_io_input_io_weiIn_bits_x_0 = PECross_165_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_181_multiply_io_input_io_weiIn_bits_last = PECross_165_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_181_multiply_io_input_io_actOut_ready = PECross_182_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_181_multiply_io_input_io_weiOut_ready = PECross_197_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_182_clock = clock;
  assign PECross_182_reset = rst;
  assign PECross_182_multiply_io_input_io_sumIn_valid = PECross_181_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_182_multiply_io_input_io_sumIn_bits_x_0 = PECross_181_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_182_multiply_io_input_io_sumIn_bits_last = PECross_181_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_182_multiply_io_input_io_sumOut_ready = PECross_183_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_182_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_182_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_182_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_182_multiply_io_input_io_actIn_valid = PECross_181_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_182_multiply_io_input_io_actIn_bits_x_0 = PECross_181_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_182_multiply_io_input_io_actIn_bits_last = PECross_181_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_182_multiply_io_input_io_weiIn_valid = PECross_166_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_182_multiply_io_input_io_weiIn_bits_x_0 = PECross_166_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_182_multiply_io_input_io_weiIn_bits_last = PECross_166_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_182_multiply_io_input_io_actOut_ready = PECross_183_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_182_multiply_io_input_io_weiOut_ready = PECross_198_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_183_clock = clock;
  assign PECross_183_reset = rst;
  assign PECross_183_multiply_io_input_io_sumIn_valid = PECross_182_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_183_multiply_io_input_io_sumIn_bits_x_0 = PECross_182_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_183_multiply_io_input_io_sumIn_bits_last = PECross_182_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_183_multiply_io_input_io_sumOut_ready = PECross_184_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_183_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_183_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_183_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_183_multiply_io_input_io_actIn_valid = PECross_182_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_183_multiply_io_input_io_actIn_bits_x_0 = PECross_182_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_183_multiply_io_input_io_actIn_bits_last = PECross_182_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_183_multiply_io_input_io_weiIn_valid = PECross_167_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_183_multiply_io_input_io_weiIn_bits_x_0 = PECross_167_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_183_multiply_io_input_io_weiIn_bits_last = PECross_167_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_183_multiply_io_input_io_actOut_ready = PECross_184_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_183_multiply_io_input_io_weiOut_ready = PECross_199_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_184_clock = clock;
  assign PECross_184_reset = rst;
  assign PECross_184_multiply_io_input_io_sumIn_valid = PECross_183_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_184_multiply_io_input_io_sumIn_bits_x_0 = PECross_183_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_184_multiply_io_input_io_sumIn_bits_last = PECross_183_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_184_multiply_io_input_io_sumOut_ready = PECross_185_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_184_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_184_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_184_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_184_multiply_io_input_io_actIn_valid = PECross_183_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_184_multiply_io_input_io_actIn_bits_x_0 = PECross_183_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_184_multiply_io_input_io_actIn_bits_last = PECross_183_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_184_multiply_io_input_io_weiIn_valid = PECross_168_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_184_multiply_io_input_io_weiIn_bits_x_0 = PECross_168_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_184_multiply_io_input_io_weiIn_bits_last = PECross_168_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_184_multiply_io_input_io_actOut_ready = PECross_185_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_184_multiply_io_input_io_weiOut_ready = PECross_200_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_185_clock = clock;
  assign PECross_185_reset = rst;
  assign PECross_185_multiply_io_input_io_sumIn_valid = PECross_184_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_185_multiply_io_input_io_sumIn_bits_x_0 = PECross_184_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_185_multiply_io_input_io_sumIn_bits_last = PECross_184_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_185_multiply_io_input_io_sumOut_ready = PECross_186_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_185_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_185_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_185_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_185_multiply_io_input_io_actIn_valid = PECross_184_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_185_multiply_io_input_io_actIn_bits_x_0 = PECross_184_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_185_multiply_io_input_io_actIn_bits_last = PECross_184_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_185_multiply_io_input_io_weiIn_valid = PECross_169_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_185_multiply_io_input_io_weiIn_bits_x_0 = PECross_169_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_185_multiply_io_input_io_weiIn_bits_last = PECross_169_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_185_multiply_io_input_io_actOut_ready = PECross_186_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_185_multiply_io_input_io_weiOut_ready = PECross_201_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_186_clock = clock;
  assign PECross_186_reset = rst;
  assign PECross_186_multiply_io_input_io_sumIn_valid = PECross_185_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_186_multiply_io_input_io_sumIn_bits_x_0 = PECross_185_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_186_multiply_io_input_io_sumIn_bits_last = PECross_185_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_186_multiply_io_input_io_sumOut_ready = PECross_187_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_186_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_186_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_186_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_186_multiply_io_input_io_actIn_valid = PECross_185_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_186_multiply_io_input_io_actIn_bits_x_0 = PECross_185_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_186_multiply_io_input_io_actIn_bits_last = PECross_185_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_186_multiply_io_input_io_weiIn_valid = PECross_170_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_186_multiply_io_input_io_weiIn_bits_x_0 = PECross_170_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_186_multiply_io_input_io_weiIn_bits_last = PECross_170_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_186_multiply_io_input_io_actOut_ready = PECross_187_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_186_multiply_io_input_io_weiOut_ready = PECross_202_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_187_clock = clock;
  assign PECross_187_reset = rst;
  assign PECross_187_multiply_io_input_io_sumIn_valid = PECross_186_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_187_multiply_io_input_io_sumIn_bits_x_0 = PECross_186_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_187_multiply_io_input_io_sumIn_bits_last = PECross_186_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_187_multiply_io_input_io_sumOut_ready = PECross_188_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_187_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_187_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_187_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_187_multiply_io_input_io_actIn_valid = PECross_186_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_187_multiply_io_input_io_actIn_bits_x_0 = PECross_186_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_187_multiply_io_input_io_actIn_bits_last = PECross_186_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_187_multiply_io_input_io_weiIn_valid = PECross_171_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_187_multiply_io_input_io_weiIn_bits_x_0 = PECross_171_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_187_multiply_io_input_io_weiIn_bits_last = PECross_171_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_187_multiply_io_input_io_actOut_ready = PECross_188_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_187_multiply_io_input_io_weiOut_ready = PECross_203_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_188_clock = clock;
  assign PECross_188_reset = rst;
  assign PECross_188_multiply_io_input_io_sumIn_valid = PECross_187_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_188_multiply_io_input_io_sumIn_bits_x_0 = PECross_187_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_188_multiply_io_input_io_sumIn_bits_last = PECross_187_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_188_multiply_io_input_io_sumOut_ready = PECross_189_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_188_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_188_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_188_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_188_multiply_io_input_io_actIn_valid = PECross_187_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_188_multiply_io_input_io_actIn_bits_x_0 = PECross_187_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_188_multiply_io_input_io_actIn_bits_last = PECross_187_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_188_multiply_io_input_io_weiIn_valid = PECross_172_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_188_multiply_io_input_io_weiIn_bits_x_0 = PECross_172_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_188_multiply_io_input_io_weiIn_bits_last = PECross_172_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_188_multiply_io_input_io_actOut_ready = PECross_189_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_188_multiply_io_input_io_weiOut_ready = PECross_204_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_189_clock = clock;
  assign PECross_189_reset = rst;
  assign PECross_189_multiply_io_input_io_sumIn_valid = PECross_188_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_189_multiply_io_input_io_sumIn_bits_x_0 = PECross_188_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_189_multiply_io_input_io_sumIn_bits_last = PECross_188_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_189_multiply_io_input_io_sumOut_ready = PECross_190_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_189_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_189_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_189_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_189_multiply_io_input_io_actIn_valid = PECross_188_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_189_multiply_io_input_io_actIn_bits_x_0 = PECross_188_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_189_multiply_io_input_io_actIn_bits_last = PECross_188_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_189_multiply_io_input_io_weiIn_valid = PECross_173_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_189_multiply_io_input_io_weiIn_bits_x_0 = PECross_173_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_189_multiply_io_input_io_weiIn_bits_last = PECross_173_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_189_multiply_io_input_io_actOut_ready = PECross_190_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_189_multiply_io_input_io_weiOut_ready = PECross_205_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_190_clock = clock;
  assign PECross_190_reset = rst;
  assign PECross_190_multiply_io_input_io_sumIn_valid = PECross_189_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_190_multiply_io_input_io_sumIn_bits_x_0 = PECross_189_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_190_multiply_io_input_io_sumIn_bits_last = PECross_189_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_190_multiply_io_input_io_sumOut_ready = PECross_191_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_190_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_190_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_190_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_190_multiply_io_input_io_actIn_valid = PECross_189_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_190_multiply_io_input_io_actIn_bits_x_0 = PECross_189_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_190_multiply_io_input_io_actIn_bits_last = PECross_189_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_190_multiply_io_input_io_weiIn_valid = PECross_174_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_190_multiply_io_input_io_weiIn_bits_x_0 = PECross_174_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_190_multiply_io_input_io_weiIn_bits_last = PECross_174_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_190_multiply_io_input_io_actOut_ready = PECross_191_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_190_multiply_io_input_io_weiOut_ready = PECross_206_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_191_clock = clock;
  assign PECross_191_reset = rst;
  assign PECross_191_multiply_io_input_io_sumIn_valid = PECross_190_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_191_multiply_io_input_io_sumIn_bits_x_0 = PECross_190_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_191_multiply_io_input_io_sumIn_bits_last = PECross_190_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_191_multiply_io_input_io_sumOut_ready = io_sumOut_11_ready; // @[mac.scala 45:29]
  assign PECross_191_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_191_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_191_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_191_multiply_io_input_io_actIn_valid = PECross_190_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_191_multiply_io_input_io_actIn_bits_x_0 = PECross_190_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_191_multiply_io_input_io_actIn_bits_last = PECross_190_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_191_multiply_io_input_io_weiIn_valid = PECross_175_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_191_multiply_io_input_io_weiIn_bits_x_0 = PECross_175_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_191_multiply_io_input_io_weiIn_bits_last = PECross_175_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_191_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_191_multiply_io_input_io_weiOut_ready = PECross_207_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_192_clock = clock;
  assign PECross_192_reset = rst;
  assign PECross_192_multiply_io_input_io_sumIn_valid = io_sumIn_12_valid; // @[mac.scala 33:28]
  assign PECross_192_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_12_bits_x_0; // @[mac.scala 33:28]
  assign PECross_192_multiply_io_input_io_sumIn_bits_last = io_sumIn_12_bits_last; // @[mac.scala 33:28]
  assign PECross_192_multiply_io_input_io_sumOut_ready = PECross_193_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_192_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_192_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_192_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_192_multiply_io_input_io_actIn_valid = io_actIn_12_valid; // @[mac.scala 32:28]
  assign PECross_192_multiply_io_input_io_actIn_bits_x_0 = io_actIn_12_bits_x_0; // @[mac.scala 32:28]
  assign PECross_192_multiply_io_input_io_actIn_bits_last = io_actIn_12_bits_last; // @[mac.scala 32:28]
  assign PECross_192_multiply_io_input_io_weiIn_valid = PECross_176_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_192_multiply_io_input_io_weiIn_bits_x_0 = PECross_176_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_192_multiply_io_input_io_weiIn_bits_last = PECross_176_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_192_multiply_io_input_io_actOut_ready = PECross_193_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_192_multiply_io_input_io_weiOut_ready = PECross_208_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_193_clock = clock;
  assign PECross_193_reset = rst;
  assign PECross_193_multiply_io_input_io_sumIn_valid = PECross_192_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_193_multiply_io_input_io_sumIn_bits_x_0 = PECross_192_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_193_multiply_io_input_io_sumIn_bits_last = PECross_192_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_193_multiply_io_input_io_sumOut_ready = PECross_194_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_193_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_193_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_193_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_193_multiply_io_input_io_actIn_valid = PECross_192_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_193_multiply_io_input_io_actIn_bits_x_0 = PECross_192_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_193_multiply_io_input_io_actIn_bits_last = PECross_192_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_193_multiply_io_input_io_weiIn_valid = PECross_177_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_193_multiply_io_input_io_weiIn_bits_x_0 = PECross_177_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_193_multiply_io_input_io_weiIn_bits_last = PECross_177_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_193_multiply_io_input_io_actOut_ready = PECross_194_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_193_multiply_io_input_io_weiOut_ready = PECross_209_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_194_clock = clock;
  assign PECross_194_reset = rst;
  assign PECross_194_multiply_io_input_io_sumIn_valid = PECross_193_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_194_multiply_io_input_io_sumIn_bits_x_0 = PECross_193_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_194_multiply_io_input_io_sumIn_bits_last = PECross_193_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_194_multiply_io_input_io_sumOut_ready = PECross_195_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_194_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_194_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_194_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_194_multiply_io_input_io_actIn_valid = PECross_193_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_194_multiply_io_input_io_actIn_bits_x_0 = PECross_193_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_194_multiply_io_input_io_actIn_bits_last = PECross_193_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_194_multiply_io_input_io_weiIn_valid = PECross_178_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_194_multiply_io_input_io_weiIn_bits_x_0 = PECross_178_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_194_multiply_io_input_io_weiIn_bits_last = PECross_178_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_194_multiply_io_input_io_actOut_ready = PECross_195_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_194_multiply_io_input_io_weiOut_ready = PECross_210_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_195_clock = clock;
  assign PECross_195_reset = rst;
  assign PECross_195_multiply_io_input_io_sumIn_valid = PECross_194_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_195_multiply_io_input_io_sumIn_bits_x_0 = PECross_194_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_195_multiply_io_input_io_sumIn_bits_last = PECross_194_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_195_multiply_io_input_io_sumOut_ready = PECross_196_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_195_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_195_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_195_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_195_multiply_io_input_io_actIn_valid = PECross_194_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_195_multiply_io_input_io_actIn_bits_x_0 = PECross_194_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_195_multiply_io_input_io_actIn_bits_last = PECross_194_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_195_multiply_io_input_io_weiIn_valid = PECross_179_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_195_multiply_io_input_io_weiIn_bits_x_0 = PECross_179_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_195_multiply_io_input_io_weiIn_bits_last = PECross_179_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_195_multiply_io_input_io_actOut_ready = PECross_196_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_195_multiply_io_input_io_weiOut_ready = PECross_211_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_196_clock = clock;
  assign PECross_196_reset = rst;
  assign PECross_196_multiply_io_input_io_sumIn_valid = PECross_195_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_196_multiply_io_input_io_sumIn_bits_x_0 = PECross_195_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_196_multiply_io_input_io_sumIn_bits_last = PECross_195_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_196_multiply_io_input_io_sumOut_ready = PECross_197_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_196_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_196_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_196_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_196_multiply_io_input_io_actIn_valid = PECross_195_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_196_multiply_io_input_io_actIn_bits_x_0 = PECross_195_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_196_multiply_io_input_io_actIn_bits_last = PECross_195_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_196_multiply_io_input_io_weiIn_valid = PECross_180_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_196_multiply_io_input_io_weiIn_bits_x_0 = PECross_180_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_196_multiply_io_input_io_weiIn_bits_last = PECross_180_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_196_multiply_io_input_io_actOut_ready = PECross_197_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_196_multiply_io_input_io_weiOut_ready = PECross_212_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_197_clock = clock;
  assign PECross_197_reset = rst;
  assign PECross_197_multiply_io_input_io_sumIn_valid = PECross_196_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_197_multiply_io_input_io_sumIn_bits_x_0 = PECross_196_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_197_multiply_io_input_io_sumIn_bits_last = PECross_196_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_197_multiply_io_input_io_sumOut_ready = PECross_198_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_197_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_197_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_197_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_197_multiply_io_input_io_actIn_valid = PECross_196_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_197_multiply_io_input_io_actIn_bits_x_0 = PECross_196_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_197_multiply_io_input_io_actIn_bits_last = PECross_196_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_197_multiply_io_input_io_weiIn_valid = PECross_181_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_197_multiply_io_input_io_weiIn_bits_x_0 = PECross_181_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_197_multiply_io_input_io_weiIn_bits_last = PECross_181_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_197_multiply_io_input_io_actOut_ready = PECross_198_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_197_multiply_io_input_io_weiOut_ready = PECross_213_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_198_clock = clock;
  assign PECross_198_reset = rst;
  assign PECross_198_multiply_io_input_io_sumIn_valid = PECross_197_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_198_multiply_io_input_io_sumIn_bits_x_0 = PECross_197_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_198_multiply_io_input_io_sumIn_bits_last = PECross_197_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_198_multiply_io_input_io_sumOut_ready = PECross_199_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_198_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_198_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_198_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_198_multiply_io_input_io_actIn_valid = PECross_197_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_198_multiply_io_input_io_actIn_bits_x_0 = PECross_197_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_198_multiply_io_input_io_actIn_bits_last = PECross_197_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_198_multiply_io_input_io_weiIn_valid = PECross_182_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_198_multiply_io_input_io_weiIn_bits_x_0 = PECross_182_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_198_multiply_io_input_io_weiIn_bits_last = PECross_182_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_198_multiply_io_input_io_actOut_ready = PECross_199_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_198_multiply_io_input_io_weiOut_ready = PECross_214_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_199_clock = clock;
  assign PECross_199_reset = rst;
  assign PECross_199_multiply_io_input_io_sumIn_valid = PECross_198_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_199_multiply_io_input_io_sumIn_bits_x_0 = PECross_198_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_199_multiply_io_input_io_sumIn_bits_last = PECross_198_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_199_multiply_io_input_io_sumOut_ready = PECross_200_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_199_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_199_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_199_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_199_multiply_io_input_io_actIn_valid = PECross_198_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_199_multiply_io_input_io_actIn_bits_x_0 = PECross_198_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_199_multiply_io_input_io_actIn_bits_last = PECross_198_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_199_multiply_io_input_io_weiIn_valid = PECross_183_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_199_multiply_io_input_io_weiIn_bits_x_0 = PECross_183_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_199_multiply_io_input_io_weiIn_bits_last = PECross_183_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_199_multiply_io_input_io_actOut_ready = PECross_200_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_199_multiply_io_input_io_weiOut_ready = PECross_215_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_200_clock = clock;
  assign PECross_200_reset = rst;
  assign PECross_200_multiply_io_input_io_sumIn_valid = PECross_199_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_200_multiply_io_input_io_sumIn_bits_x_0 = PECross_199_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_200_multiply_io_input_io_sumIn_bits_last = PECross_199_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_200_multiply_io_input_io_sumOut_ready = PECross_201_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_200_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_200_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_200_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_200_multiply_io_input_io_actIn_valid = PECross_199_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_200_multiply_io_input_io_actIn_bits_x_0 = PECross_199_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_200_multiply_io_input_io_actIn_bits_last = PECross_199_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_200_multiply_io_input_io_weiIn_valid = PECross_184_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_200_multiply_io_input_io_weiIn_bits_x_0 = PECross_184_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_200_multiply_io_input_io_weiIn_bits_last = PECross_184_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_200_multiply_io_input_io_actOut_ready = PECross_201_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_200_multiply_io_input_io_weiOut_ready = PECross_216_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_201_clock = clock;
  assign PECross_201_reset = rst;
  assign PECross_201_multiply_io_input_io_sumIn_valid = PECross_200_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_201_multiply_io_input_io_sumIn_bits_x_0 = PECross_200_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_201_multiply_io_input_io_sumIn_bits_last = PECross_200_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_201_multiply_io_input_io_sumOut_ready = PECross_202_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_201_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_201_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_201_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_201_multiply_io_input_io_actIn_valid = PECross_200_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_201_multiply_io_input_io_actIn_bits_x_0 = PECross_200_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_201_multiply_io_input_io_actIn_bits_last = PECross_200_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_201_multiply_io_input_io_weiIn_valid = PECross_185_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_201_multiply_io_input_io_weiIn_bits_x_0 = PECross_185_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_201_multiply_io_input_io_weiIn_bits_last = PECross_185_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_201_multiply_io_input_io_actOut_ready = PECross_202_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_201_multiply_io_input_io_weiOut_ready = PECross_217_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_202_clock = clock;
  assign PECross_202_reset = rst;
  assign PECross_202_multiply_io_input_io_sumIn_valid = PECross_201_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_202_multiply_io_input_io_sumIn_bits_x_0 = PECross_201_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_202_multiply_io_input_io_sumIn_bits_last = PECross_201_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_202_multiply_io_input_io_sumOut_ready = PECross_203_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_202_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_202_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_202_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_202_multiply_io_input_io_actIn_valid = PECross_201_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_202_multiply_io_input_io_actIn_bits_x_0 = PECross_201_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_202_multiply_io_input_io_actIn_bits_last = PECross_201_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_202_multiply_io_input_io_weiIn_valid = PECross_186_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_202_multiply_io_input_io_weiIn_bits_x_0 = PECross_186_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_202_multiply_io_input_io_weiIn_bits_last = PECross_186_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_202_multiply_io_input_io_actOut_ready = PECross_203_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_202_multiply_io_input_io_weiOut_ready = PECross_218_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_203_clock = clock;
  assign PECross_203_reset = rst;
  assign PECross_203_multiply_io_input_io_sumIn_valid = PECross_202_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_203_multiply_io_input_io_sumIn_bits_x_0 = PECross_202_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_203_multiply_io_input_io_sumIn_bits_last = PECross_202_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_203_multiply_io_input_io_sumOut_ready = PECross_204_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_203_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_203_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_203_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_203_multiply_io_input_io_actIn_valid = PECross_202_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_203_multiply_io_input_io_actIn_bits_x_0 = PECross_202_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_203_multiply_io_input_io_actIn_bits_last = PECross_202_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_203_multiply_io_input_io_weiIn_valid = PECross_187_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_203_multiply_io_input_io_weiIn_bits_x_0 = PECross_187_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_203_multiply_io_input_io_weiIn_bits_last = PECross_187_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_203_multiply_io_input_io_actOut_ready = PECross_204_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_203_multiply_io_input_io_weiOut_ready = PECross_219_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_204_clock = clock;
  assign PECross_204_reset = rst;
  assign PECross_204_multiply_io_input_io_sumIn_valid = PECross_203_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_204_multiply_io_input_io_sumIn_bits_x_0 = PECross_203_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_204_multiply_io_input_io_sumIn_bits_last = PECross_203_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_204_multiply_io_input_io_sumOut_ready = PECross_205_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_204_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_204_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_204_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_204_multiply_io_input_io_actIn_valid = PECross_203_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_204_multiply_io_input_io_actIn_bits_x_0 = PECross_203_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_204_multiply_io_input_io_actIn_bits_last = PECross_203_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_204_multiply_io_input_io_weiIn_valid = PECross_188_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_204_multiply_io_input_io_weiIn_bits_x_0 = PECross_188_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_204_multiply_io_input_io_weiIn_bits_last = PECross_188_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_204_multiply_io_input_io_actOut_ready = PECross_205_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_204_multiply_io_input_io_weiOut_ready = PECross_220_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_205_clock = clock;
  assign PECross_205_reset = rst;
  assign PECross_205_multiply_io_input_io_sumIn_valid = PECross_204_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_205_multiply_io_input_io_sumIn_bits_x_0 = PECross_204_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_205_multiply_io_input_io_sumIn_bits_last = PECross_204_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_205_multiply_io_input_io_sumOut_ready = PECross_206_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_205_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_205_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_205_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_205_multiply_io_input_io_actIn_valid = PECross_204_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_205_multiply_io_input_io_actIn_bits_x_0 = PECross_204_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_205_multiply_io_input_io_actIn_bits_last = PECross_204_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_205_multiply_io_input_io_weiIn_valid = PECross_189_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_205_multiply_io_input_io_weiIn_bits_x_0 = PECross_189_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_205_multiply_io_input_io_weiIn_bits_last = PECross_189_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_205_multiply_io_input_io_actOut_ready = PECross_206_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_205_multiply_io_input_io_weiOut_ready = PECross_221_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_206_clock = clock;
  assign PECross_206_reset = rst;
  assign PECross_206_multiply_io_input_io_sumIn_valid = PECross_205_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_206_multiply_io_input_io_sumIn_bits_x_0 = PECross_205_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_206_multiply_io_input_io_sumIn_bits_last = PECross_205_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_206_multiply_io_input_io_sumOut_ready = PECross_207_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_206_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_206_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_206_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_206_multiply_io_input_io_actIn_valid = PECross_205_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_206_multiply_io_input_io_actIn_bits_x_0 = PECross_205_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_206_multiply_io_input_io_actIn_bits_last = PECross_205_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_206_multiply_io_input_io_weiIn_valid = PECross_190_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_206_multiply_io_input_io_weiIn_bits_x_0 = PECross_190_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_206_multiply_io_input_io_weiIn_bits_last = PECross_190_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_206_multiply_io_input_io_actOut_ready = PECross_207_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_206_multiply_io_input_io_weiOut_ready = PECross_222_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_207_clock = clock;
  assign PECross_207_reset = rst;
  assign PECross_207_multiply_io_input_io_sumIn_valid = PECross_206_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_207_multiply_io_input_io_sumIn_bits_x_0 = PECross_206_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_207_multiply_io_input_io_sumIn_bits_last = PECross_206_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_207_multiply_io_input_io_sumOut_ready = io_sumOut_12_ready; // @[mac.scala 45:29]
  assign PECross_207_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_207_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_207_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_207_multiply_io_input_io_actIn_valid = PECross_206_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_207_multiply_io_input_io_actIn_bits_x_0 = PECross_206_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_207_multiply_io_input_io_actIn_bits_last = PECross_206_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_207_multiply_io_input_io_weiIn_valid = PECross_191_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_207_multiply_io_input_io_weiIn_bits_x_0 = PECross_191_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_207_multiply_io_input_io_weiIn_bits_last = PECross_191_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_207_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_207_multiply_io_input_io_weiOut_ready = PECross_223_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_208_clock = clock;
  assign PECross_208_reset = rst;
  assign PECross_208_multiply_io_input_io_sumIn_valid = io_sumIn_13_valid; // @[mac.scala 33:28]
  assign PECross_208_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_13_bits_x_0; // @[mac.scala 33:28]
  assign PECross_208_multiply_io_input_io_sumIn_bits_last = io_sumIn_13_bits_last; // @[mac.scala 33:28]
  assign PECross_208_multiply_io_input_io_sumOut_ready = PECross_209_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_208_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_208_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_208_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_208_multiply_io_input_io_actIn_valid = io_actIn_13_valid; // @[mac.scala 32:28]
  assign PECross_208_multiply_io_input_io_actIn_bits_x_0 = io_actIn_13_bits_x_0; // @[mac.scala 32:28]
  assign PECross_208_multiply_io_input_io_actIn_bits_last = io_actIn_13_bits_last; // @[mac.scala 32:28]
  assign PECross_208_multiply_io_input_io_weiIn_valid = PECross_192_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_208_multiply_io_input_io_weiIn_bits_x_0 = PECross_192_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_208_multiply_io_input_io_weiIn_bits_last = PECross_192_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_208_multiply_io_input_io_actOut_ready = PECross_209_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_208_multiply_io_input_io_weiOut_ready = PECross_224_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_209_clock = clock;
  assign PECross_209_reset = rst;
  assign PECross_209_multiply_io_input_io_sumIn_valid = PECross_208_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_209_multiply_io_input_io_sumIn_bits_x_0 = PECross_208_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_209_multiply_io_input_io_sumIn_bits_last = PECross_208_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_209_multiply_io_input_io_sumOut_ready = PECross_210_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_209_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_209_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_209_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_209_multiply_io_input_io_actIn_valid = PECross_208_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_209_multiply_io_input_io_actIn_bits_x_0 = PECross_208_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_209_multiply_io_input_io_actIn_bits_last = PECross_208_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_209_multiply_io_input_io_weiIn_valid = PECross_193_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_209_multiply_io_input_io_weiIn_bits_x_0 = PECross_193_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_209_multiply_io_input_io_weiIn_bits_last = PECross_193_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_209_multiply_io_input_io_actOut_ready = PECross_210_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_209_multiply_io_input_io_weiOut_ready = PECross_225_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_210_clock = clock;
  assign PECross_210_reset = rst;
  assign PECross_210_multiply_io_input_io_sumIn_valid = PECross_209_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_210_multiply_io_input_io_sumIn_bits_x_0 = PECross_209_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_210_multiply_io_input_io_sumIn_bits_last = PECross_209_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_210_multiply_io_input_io_sumOut_ready = PECross_211_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_210_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_210_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_210_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_210_multiply_io_input_io_actIn_valid = PECross_209_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_210_multiply_io_input_io_actIn_bits_x_0 = PECross_209_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_210_multiply_io_input_io_actIn_bits_last = PECross_209_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_210_multiply_io_input_io_weiIn_valid = PECross_194_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_210_multiply_io_input_io_weiIn_bits_x_0 = PECross_194_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_210_multiply_io_input_io_weiIn_bits_last = PECross_194_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_210_multiply_io_input_io_actOut_ready = PECross_211_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_210_multiply_io_input_io_weiOut_ready = PECross_226_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_211_clock = clock;
  assign PECross_211_reset = rst;
  assign PECross_211_multiply_io_input_io_sumIn_valid = PECross_210_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_211_multiply_io_input_io_sumIn_bits_x_0 = PECross_210_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_211_multiply_io_input_io_sumIn_bits_last = PECross_210_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_211_multiply_io_input_io_sumOut_ready = PECross_212_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_211_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_211_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_211_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_211_multiply_io_input_io_actIn_valid = PECross_210_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_211_multiply_io_input_io_actIn_bits_x_0 = PECross_210_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_211_multiply_io_input_io_actIn_bits_last = PECross_210_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_211_multiply_io_input_io_weiIn_valid = PECross_195_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_211_multiply_io_input_io_weiIn_bits_x_0 = PECross_195_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_211_multiply_io_input_io_weiIn_bits_last = PECross_195_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_211_multiply_io_input_io_actOut_ready = PECross_212_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_211_multiply_io_input_io_weiOut_ready = PECross_227_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_212_clock = clock;
  assign PECross_212_reset = rst;
  assign PECross_212_multiply_io_input_io_sumIn_valid = PECross_211_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_212_multiply_io_input_io_sumIn_bits_x_0 = PECross_211_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_212_multiply_io_input_io_sumIn_bits_last = PECross_211_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_212_multiply_io_input_io_sumOut_ready = PECross_213_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_212_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_212_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_212_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_212_multiply_io_input_io_actIn_valid = PECross_211_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_212_multiply_io_input_io_actIn_bits_x_0 = PECross_211_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_212_multiply_io_input_io_actIn_bits_last = PECross_211_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_212_multiply_io_input_io_weiIn_valid = PECross_196_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_212_multiply_io_input_io_weiIn_bits_x_0 = PECross_196_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_212_multiply_io_input_io_weiIn_bits_last = PECross_196_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_212_multiply_io_input_io_actOut_ready = PECross_213_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_212_multiply_io_input_io_weiOut_ready = PECross_228_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_213_clock = clock;
  assign PECross_213_reset = rst;
  assign PECross_213_multiply_io_input_io_sumIn_valid = PECross_212_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_213_multiply_io_input_io_sumIn_bits_x_0 = PECross_212_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_213_multiply_io_input_io_sumIn_bits_last = PECross_212_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_213_multiply_io_input_io_sumOut_ready = PECross_214_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_213_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_213_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_213_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_213_multiply_io_input_io_actIn_valid = PECross_212_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_213_multiply_io_input_io_actIn_bits_x_0 = PECross_212_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_213_multiply_io_input_io_actIn_bits_last = PECross_212_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_213_multiply_io_input_io_weiIn_valid = PECross_197_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_213_multiply_io_input_io_weiIn_bits_x_0 = PECross_197_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_213_multiply_io_input_io_weiIn_bits_last = PECross_197_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_213_multiply_io_input_io_actOut_ready = PECross_214_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_213_multiply_io_input_io_weiOut_ready = PECross_229_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_214_clock = clock;
  assign PECross_214_reset = rst;
  assign PECross_214_multiply_io_input_io_sumIn_valid = PECross_213_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_214_multiply_io_input_io_sumIn_bits_x_0 = PECross_213_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_214_multiply_io_input_io_sumIn_bits_last = PECross_213_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_214_multiply_io_input_io_sumOut_ready = PECross_215_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_214_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_214_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_214_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_214_multiply_io_input_io_actIn_valid = PECross_213_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_214_multiply_io_input_io_actIn_bits_x_0 = PECross_213_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_214_multiply_io_input_io_actIn_bits_last = PECross_213_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_214_multiply_io_input_io_weiIn_valid = PECross_198_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_214_multiply_io_input_io_weiIn_bits_x_0 = PECross_198_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_214_multiply_io_input_io_weiIn_bits_last = PECross_198_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_214_multiply_io_input_io_actOut_ready = PECross_215_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_214_multiply_io_input_io_weiOut_ready = PECross_230_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_215_clock = clock;
  assign PECross_215_reset = rst;
  assign PECross_215_multiply_io_input_io_sumIn_valid = PECross_214_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_215_multiply_io_input_io_sumIn_bits_x_0 = PECross_214_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_215_multiply_io_input_io_sumIn_bits_last = PECross_214_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_215_multiply_io_input_io_sumOut_ready = PECross_216_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_215_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_215_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_215_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_215_multiply_io_input_io_actIn_valid = PECross_214_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_215_multiply_io_input_io_actIn_bits_x_0 = PECross_214_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_215_multiply_io_input_io_actIn_bits_last = PECross_214_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_215_multiply_io_input_io_weiIn_valid = PECross_199_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_215_multiply_io_input_io_weiIn_bits_x_0 = PECross_199_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_215_multiply_io_input_io_weiIn_bits_last = PECross_199_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_215_multiply_io_input_io_actOut_ready = PECross_216_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_215_multiply_io_input_io_weiOut_ready = PECross_231_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_216_clock = clock;
  assign PECross_216_reset = rst;
  assign PECross_216_multiply_io_input_io_sumIn_valid = PECross_215_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_216_multiply_io_input_io_sumIn_bits_x_0 = PECross_215_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_216_multiply_io_input_io_sumIn_bits_last = PECross_215_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_216_multiply_io_input_io_sumOut_ready = PECross_217_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_216_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_216_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_216_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_216_multiply_io_input_io_actIn_valid = PECross_215_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_216_multiply_io_input_io_actIn_bits_x_0 = PECross_215_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_216_multiply_io_input_io_actIn_bits_last = PECross_215_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_216_multiply_io_input_io_weiIn_valid = PECross_200_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_216_multiply_io_input_io_weiIn_bits_x_0 = PECross_200_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_216_multiply_io_input_io_weiIn_bits_last = PECross_200_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_216_multiply_io_input_io_actOut_ready = PECross_217_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_216_multiply_io_input_io_weiOut_ready = PECross_232_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_217_clock = clock;
  assign PECross_217_reset = rst;
  assign PECross_217_multiply_io_input_io_sumIn_valid = PECross_216_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_217_multiply_io_input_io_sumIn_bits_x_0 = PECross_216_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_217_multiply_io_input_io_sumIn_bits_last = PECross_216_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_217_multiply_io_input_io_sumOut_ready = PECross_218_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_217_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_217_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_217_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_217_multiply_io_input_io_actIn_valid = PECross_216_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_217_multiply_io_input_io_actIn_bits_x_0 = PECross_216_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_217_multiply_io_input_io_actIn_bits_last = PECross_216_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_217_multiply_io_input_io_weiIn_valid = PECross_201_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_217_multiply_io_input_io_weiIn_bits_x_0 = PECross_201_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_217_multiply_io_input_io_weiIn_bits_last = PECross_201_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_217_multiply_io_input_io_actOut_ready = PECross_218_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_217_multiply_io_input_io_weiOut_ready = PECross_233_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_218_clock = clock;
  assign PECross_218_reset = rst;
  assign PECross_218_multiply_io_input_io_sumIn_valid = PECross_217_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_218_multiply_io_input_io_sumIn_bits_x_0 = PECross_217_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_218_multiply_io_input_io_sumIn_bits_last = PECross_217_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_218_multiply_io_input_io_sumOut_ready = PECross_219_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_218_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_218_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_218_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_218_multiply_io_input_io_actIn_valid = PECross_217_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_218_multiply_io_input_io_actIn_bits_x_0 = PECross_217_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_218_multiply_io_input_io_actIn_bits_last = PECross_217_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_218_multiply_io_input_io_weiIn_valid = PECross_202_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_218_multiply_io_input_io_weiIn_bits_x_0 = PECross_202_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_218_multiply_io_input_io_weiIn_bits_last = PECross_202_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_218_multiply_io_input_io_actOut_ready = PECross_219_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_218_multiply_io_input_io_weiOut_ready = PECross_234_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_219_clock = clock;
  assign PECross_219_reset = rst;
  assign PECross_219_multiply_io_input_io_sumIn_valid = PECross_218_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_219_multiply_io_input_io_sumIn_bits_x_0 = PECross_218_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_219_multiply_io_input_io_sumIn_bits_last = PECross_218_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_219_multiply_io_input_io_sumOut_ready = PECross_220_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_219_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_219_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_219_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_219_multiply_io_input_io_actIn_valid = PECross_218_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_219_multiply_io_input_io_actIn_bits_x_0 = PECross_218_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_219_multiply_io_input_io_actIn_bits_last = PECross_218_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_219_multiply_io_input_io_weiIn_valid = PECross_203_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_219_multiply_io_input_io_weiIn_bits_x_0 = PECross_203_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_219_multiply_io_input_io_weiIn_bits_last = PECross_203_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_219_multiply_io_input_io_actOut_ready = PECross_220_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_219_multiply_io_input_io_weiOut_ready = PECross_235_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_220_clock = clock;
  assign PECross_220_reset = rst;
  assign PECross_220_multiply_io_input_io_sumIn_valid = PECross_219_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_220_multiply_io_input_io_sumIn_bits_x_0 = PECross_219_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_220_multiply_io_input_io_sumIn_bits_last = PECross_219_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_220_multiply_io_input_io_sumOut_ready = PECross_221_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_220_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_220_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_220_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_220_multiply_io_input_io_actIn_valid = PECross_219_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_220_multiply_io_input_io_actIn_bits_x_0 = PECross_219_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_220_multiply_io_input_io_actIn_bits_last = PECross_219_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_220_multiply_io_input_io_weiIn_valid = PECross_204_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_220_multiply_io_input_io_weiIn_bits_x_0 = PECross_204_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_220_multiply_io_input_io_weiIn_bits_last = PECross_204_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_220_multiply_io_input_io_actOut_ready = PECross_221_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_220_multiply_io_input_io_weiOut_ready = PECross_236_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_221_clock = clock;
  assign PECross_221_reset = rst;
  assign PECross_221_multiply_io_input_io_sumIn_valid = PECross_220_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_221_multiply_io_input_io_sumIn_bits_x_0 = PECross_220_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_221_multiply_io_input_io_sumIn_bits_last = PECross_220_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_221_multiply_io_input_io_sumOut_ready = PECross_222_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_221_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_221_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_221_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_221_multiply_io_input_io_actIn_valid = PECross_220_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_221_multiply_io_input_io_actIn_bits_x_0 = PECross_220_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_221_multiply_io_input_io_actIn_bits_last = PECross_220_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_221_multiply_io_input_io_weiIn_valid = PECross_205_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_221_multiply_io_input_io_weiIn_bits_x_0 = PECross_205_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_221_multiply_io_input_io_weiIn_bits_last = PECross_205_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_221_multiply_io_input_io_actOut_ready = PECross_222_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_221_multiply_io_input_io_weiOut_ready = PECross_237_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_222_clock = clock;
  assign PECross_222_reset = rst;
  assign PECross_222_multiply_io_input_io_sumIn_valid = PECross_221_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_222_multiply_io_input_io_sumIn_bits_x_0 = PECross_221_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_222_multiply_io_input_io_sumIn_bits_last = PECross_221_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_222_multiply_io_input_io_sumOut_ready = PECross_223_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_222_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_222_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_222_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_222_multiply_io_input_io_actIn_valid = PECross_221_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_222_multiply_io_input_io_actIn_bits_x_0 = PECross_221_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_222_multiply_io_input_io_actIn_bits_last = PECross_221_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_222_multiply_io_input_io_weiIn_valid = PECross_206_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_222_multiply_io_input_io_weiIn_bits_x_0 = PECross_206_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_222_multiply_io_input_io_weiIn_bits_last = PECross_206_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_222_multiply_io_input_io_actOut_ready = PECross_223_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_222_multiply_io_input_io_weiOut_ready = PECross_238_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_223_clock = clock;
  assign PECross_223_reset = rst;
  assign PECross_223_multiply_io_input_io_sumIn_valid = PECross_222_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_223_multiply_io_input_io_sumIn_bits_x_0 = PECross_222_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_223_multiply_io_input_io_sumIn_bits_last = PECross_222_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_223_multiply_io_input_io_sumOut_ready = io_sumOut_13_ready; // @[mac.scala 45:29]
  assign PECross_223_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_223_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_223_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_223_multiply_io_input_io_actIn_valid = PECross_222_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_223_multiply_io_input_io_actIn_bits_x_0 = PECross_222_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_223_multiply_io_input_io_actIn_bits_last = PECross_222_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_223_multiply_io_input_io_weiIn_valid = PECross_207_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_223_multiply_io_input_io_weiIn_bits_x_0 = PECross_207_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_223_multiply_io_input_io_weiIn_bits_last = PECross_207_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_223_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_223_multiply_io_input_io_weiOut_ready = PECross_239_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_224_clock = clock;
  assign PECross_224_reset = rst;
  assign PECross_224_multiply_io_input_io_sumIn_valid = io_sumIn_14_valid; // @[mac.scala 33:28]
  assign PECross_224_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_14_bits_x_0; // @[mac.scala 33:28]
  assign PECross_224_multiply_io_input_io_sumIn_bits_last = io_sumIn_14_bits_last; // @[mac.scala 33:28]
  assign PECross_224_multiply_io_input_io_sumOut_ready = PECross_225_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_224_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_224_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_224_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_224_multiply_io_input_io_actIn_valid = io_actIn_14_valid; // @[mac.scala 32:28]
  assign PECross_224_multiply_io_input_io_actIn_bits_x_0 = io_actIn_14_bits_x_0; // @[mac.scala 32:28]
  assign PECross_224_multiply_io_input_io_actIn_bits_last = io_actIn_14_bits_last; // @[mac.scala 32:28]
  assign PECross_224_multiply_io_input_io_weiIn_valid = PECross_208_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_224_multiply_io_input_io_weiIn_bits_x_0 = PECross_208_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_224_multiply_io_input_io_weiIn_bits_last = PECross_208_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_224_multiply_io_input_io_actOut_ready = PECross_225_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_224_multiply_io_input_io_weiOut_ready = PECross_240_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_225_clock = clock;
  assign PECross_225_reset = rst;
  assign PECross_225_multiply_io_input_io_sumIn_valid = PECross_224_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_225_multiply_io_input_io_sumIn_bits_x_0 = PECross_224_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_225_multiply_io_input_io_sumIn_bits_last = PECross_224_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_225_multiply_io_input_io_sumOut_ready = PECross_226_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_225_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_225_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_225_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_225_multiply_io_input_io_actIn_valid = PECross_224_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_225_multiply_io_input_io_actIn_bits_x_0 = PECross_224_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_225_multiply_io_input_io_actIn_bits_last = PECross_224_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_225_multiply_io_input_io_weiIn_valid = PECross_209_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_225_multiply_io_input_io_weiIn_bits_x_0 = PECross_209_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_225_multiply_io_input_io_weiIn_bits_last = PECross_209_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_225_multiply_io_input_io_actOut_ready = PECross_226_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_225_multiply_io_input_io_weiOut_ready = PECross_241_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_226_clock = clock;
  assign PECross_226_reset = rst;
  assign PECross_226_multiply_io_input_io_sumIn_valid = PECross_225_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_226_multiply_io_input_io_sumIn_bits_x_0 = PECross_225_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_226_multiply_io_input_io_sumIn_bits_last = PECross_225_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_226_multiply_io_input_io_sumOut_ready = PECross_227_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_226_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_226_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_226_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_226_multiply_io_input_io_actIn_valid = PECross_225_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_226_multiply_io_input_io_actIn_bits_x_0 = PECross_225_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_226_multiply_io_input_io_actIn_bits_last = PECross_225_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_226_multiply_io_input_io_weiIn_valid = PECross_210_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_226_multiply_io_input_io_weiIn_bits_x_0 = PECross_210_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_226_multiply_io_input_io_weiIn_bits_last = PECross_210_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_226_multiply_io_input_io_actOut_ready = PECross_227_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_226_multiply_io_input_io_weiOut_ready = PECross_242_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_227_clock = clock;
  assign PECross_227_reset = rst;
  assign PECross_227_multiply_io_input_io_sumIn_valid = PECross_226_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_227_multiply_io_input_io_sumIn_bits_x_0 = PECross_226_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_227_multiply_io_input_io_sumIn_bits_last = PECross_226_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_227_multiply_io_input_io_sumOut_ready = PECross_228_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_227_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_227_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_227_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_227_multiply_io_input_io_actIn_valid = PECross_226_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_227_multiply_io_input_io_actIn_bits_x_0 = PECross_226_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_227_multiply_io_input_io_actIn_bits_last = PECross_226_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_227_multiply_io_input_io_weiIn_valid = PECross_211_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_227_multiply_io_input_io_weiIn_bits_x_0 = PECross_211_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_227_multiply_io_input_io_weiIn_bits_last = PECross_211_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_227_multiply_io_input_io_actOut_ready = PECross_228_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_227_multiply_io_input_io_weiOut_ready = PECross_243_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_228_clock = clock;
  assign PECross_228_reset = rst;
  assign PECross_228_multiply_io_input_io_sumIn_valid = PECross_227_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_228_multiply_io_input_io_sumIn_bits_x_0 = PECross_227_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_228_multiply_io_input_io_sumIn_bits_last = PECross_227_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_228_multiply_io_input_io_sumOut_ready = PECross_229_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_228_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_228_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_228_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_228_multiply_io_input_io_actIn_valid = PECross_227_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_228_multiply_io_input_io_actIn_bits_x_0 = PECross_227_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_228_multiply_io_input_io_actIn_bits_last = PECross_227_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_228_multiply_io_input_io_weiIn_valid = PECross_212_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_228_multiply_io_input_io_weiIn_bits_x_0 = PECross_212_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_228_multiply_io_input_io_weiIn_bits_last = PECross_212_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_228_multiply_io_input_io_actOut_ready = PECross_229_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_228_multiply_io_input_io_weiOut_ready = PECross_244_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_229_clock = clock;
  assign PECross_229_reset = rst;
  assign PECross_229_multiply_io_input_io_sumIn_valid = PECross_228_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_229_multiply_io_input_io_sumIn_bits_x_0 = PECross_228_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_229_multiply_io_input_io_sumIn_bits_last = PECross_228_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_229_multiply_io_input_io_sumOut_ready = PECross_230_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_229_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_229_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_229_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_229_multiply_io_input_io_actIn_valid = PECross_228_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_229_multiply_io_input_io_actIn_bits_x_0 = PECross_228_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_229_multiply_io_input_io_actIn_bits_last = PECross_228_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_229_multiply_io_input_io_weiIn_valid = PECross_213_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_229_multiply_io_input_io_weiIn_bits_x_0 = PECross_213_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_229_multiply_io_input_io_weiIn_bits_last = PECross_213_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_229_multiply_io_input_io_actOut_ready = PECross_230_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_229_multiply_io_input_io_weiOut_ready = PECross_245_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_230_clock = clock;
  assign PECross_230_reset = rst;
  assign PECross_230_multiply_io_input_io_sumIn_valid = PECross_229_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_230_multiply_io_input_io_sumIn_bits_x_0 = PECross_229_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_230_multiply_io_input_io_sumIn_bits_last = PECross_229_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_230_multiply_io_input_io_sumOut_ready = PECross_231_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_230_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_230_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_230_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_230_multiply_io_input_io_actIn_valid = PECross_229_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_230_multiply_io_input_io_actIn_bits_x_0 = PECross_229_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_230_multiply_io_input_io_actIn_bits_last = PECross_229_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_230_multiply_io_input_io_weiIn_valid = PECross_214_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_230_multiply_io_input_io_weiIn_bits_x_0 = PECross_214_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_230_multiply_io_input_io_weiIn_bits_last = PECross_214_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_230_multiply_io_input_io_actOut_ready = PECross_231_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_230_multiply_io_input_io_weiOut_ready = PECross_246_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_231_clock = clock;
  assign PECross_231_reset = rst;
  assign PECross_231_multiply_io_input_io_sumIn_valid = PECross_230_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_231_multiply_io_input_io_sumIn_bits_x_0 = PECross_230_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_231_multiply_io_input_io_sumIn_bits_last = PECross_230_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_231_multiply_io_input_io_sumOut_ready = PECross_232_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_231_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_231_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_231_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_231_multiply_io_input_io_actIn_valid = PECross_230_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_231_multiply_io_input_io_actIn_bits_x_0 = PECross_230_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_231_multiply_io_input_io_actIn_bits_last = PECross_230_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_231_multiply_io_input_io_weiIn_valid = PECross_215_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_231_multiply_io_input_io_weiIn_bits_x_0 = PECross_215_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_231_multiply_io_input_io_weiIn_bits_last = PECross_215_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_231_multiply_io_input_io_actOut_ready = PECross_232_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_231_multiply_io_input_io_weiOut_ready = PECross_247_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_232_clock = clock;
  assign PECross_232_reset = rst;
  assign PECross_232_multiply_io_input_io_sumIn_valid = PECross_231_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_232_multiply_io_input_io_sumIn_bits_x_0 = PECross_231_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_232_multiply_io_input_io_sumIn_bits_last = PECross_231_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_232_multiply_io_input_io_sumOut_ready = PECross_233_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_232_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_232_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_232_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_232_multiply_io_input_io_actIn_valid = PECross_231_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_232_multiply_io_input_io_actIn_bits_x_0 = PECross_231_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_232_multiply_io_input_io_actIn_bits_last = PECross_231_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_232_multiply_io_input_io_weiIn_valid = PECross_216_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_232_multiply_io_input_io_weiIn_bits_x_0 = PECross_216_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_232_multiply_io_input_io_weiIn_bits_last = PECross_216_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_232_multiply_io_input_io_actOut_ready = PECross_233_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_232_multiply_io_input_io_weiOut_ready = PECross_248_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_233_clock = clock;
  assign PECross_233_reset = rst;
  assign PECross_233_multiply_io_input_io_sumIn_valid = PECross_232_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_233_multiply_io_input_io_sumIn_bits_x_0 = PECross_232_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_233_multiply_io_input_io_sumIn_bits_last = PECross_232_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_233_multiply_io_input_io_sumOut_ready = PECross_234_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_233_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_233_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_233_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_233_multiply_io_input_io_actIn_valid = PECross_232_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_233_multiply_io_input_io_actIn_bits_x_0 = PECross_232_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_233_multiply_io_input_io_actIn_bits_last = PECross_232_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_233_multiply_io_input_io_weiIn_valid = PECross_217_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_233_multiply_io_input_io_weiIn_bits_x_0 = PECross_217_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_233_multiply_io_input_io_weiIn_bits_last = PECross_217_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_233_multiply_io_input_io_actOut_ready = PECross_234_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_233_multiply_io_input_io_weiOut_ready = PECross_249_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_234_clock = clock;
  assign PECross_234_reset = rst;
  assign PECross_234_multiply_io_input_io_sumIn_valid = PECross_233_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_234_multiply_io_input_io_sumIn_bits_x_0 = PECross_233_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_234_multiply_io_input_io_sumIn_bits_last = PECross_233_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_234_multiply_io_input_io_sumOut_ready = PECross_235_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_234_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_234_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_234_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_234_multiply_io_input_io_actIn_valid = PECross_233_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_234_multiply_io_input_io_actIn_bits_x_0 = PECross_233_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_234_multiply_io_input_io_actIn_bits_last = PECross_233_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_234_multiply_io_input_io_weiIn_valid = PECross_218_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_234_multiply_io_input_io_weiIn_bits_x_0 = PECross_218_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_234_multiply_io_input_io_weiIn_bits_last = PECross_218_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_234_multiply_io_input_io_actOut_ready = PECross_235_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_234_multiply_io_input_io_weiOut_ready = PECross_250_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_235_clock = clock;
  assign PECross_235_reset = rst;
  assign PECross_235_multiply_io_input_io_sumIn_valid = PECross_234_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_235_multiply_io_input_io_sumIn_bits_x_0 = PECross_234_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_235_multiply_io_input_io_sumIn_bits_last = PECross_234_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_235_multiply_io_input_io_sumOut_ready = PECross_236_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_235_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_235_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_235_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_235_multiply_io_input_io_actIn_valid = PECross_234_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_235_multiply_io_input_io_actIn_bits_x_0 = PECross_234_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_235_multiply_io_input_io_actIn_bits_last = PECross_234_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_235_multiply_io_input_io_weiIn_valid = PECross_219_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_235_multiply_io_input_io_weiIn_bits_x_0 = PECross_219_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_235_multiply_io_input_io_weiIn_bits_last = PECross_219_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_235_multiply_io_input_io_actOut_ready = PECross_236_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_235_multiply_io_input_io_weiOut_ready = PECross_251_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_236_clock = clock;
  assign PECross_236_reset = rst;
  assign PECross_236_multiply_io_input_io_sumIn_valid = PECross_235_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_236_multiply_io_input_io_sumIn_bits_x_0 = PECross_235_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_236_multiply_io_input_io_sumIn_bits_last = PECross_235_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_236_multiply_io_input_io_sumOut_ready = PECross_237_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_236_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_236_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_236_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_236_multiply_io_input_io_actIn_valid = PECross_235_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_236_multiply_io_input_io_actIn_bits_x_0 = PECross_235_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_236_multiply_io_input_io_actIn_bits_last = PECross_235_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_236_multiply_io_input_io_weiIn_valid = PECross_220_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_236_multiply_io_input_io_weiIn_bits_x_0 = PECross_220_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_236_multiply_io_input_io_weiIn_bits_last = PECross_220_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_236_multiply_io_input_io_actOut_ready = PECross_237_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_236_multiply_io_input_io_weiOut_ready = PECross_252_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_237_clock = clock;
  assign PECross_237_reset = rst;
  assign PECross_237_multiply_io_input_io_sumIn_valid = PECross_236_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_237_multiply_io_input_io_sumIn_bits_x_0 = PECross_236_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_237_multiply_io_input_io_sumIn_bits_last = PECross_236_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_237_multiply_io_input_io_sumOut_ready = PECross_238_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_237_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_237_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_237_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_237_multiply_io_input_io_actIn_valid = PECross_236_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_237_multiply_io_input_io_actIn_bits_x_0 = PECross_236_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_237_multiply_io_input_io_actIn_bits_last = PECross_236_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_237_multiply_io_input_io_weiIn_valid = PECross_221_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_237_multiply_io_input_io_weiIn_bits_x_0 = PECross_221_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_237_multiply_io_input_io_weiIn_bits_last = PECross_221_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_237_multiply_io_input_io_actOut_ready = PECross_238_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_237_multiply_io_input_io_weiOut_ready = PECross_253_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_238_clock = clock;
  assign PECross_238_reset = rst;
  assign PECross_238_multiply_io_input_io_sumIn_valid = PECross_237_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_238_multiply_io_input_io_sumIn_bits_x_0 = PECross_237_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_238_multiply_io_input_io_sumIn_bits_last = PECross_237_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_238_multiply_io_input_io_sumOut_ready = PECross_239_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_238_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_238_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_238_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_238_multiply_io_input_io_actIn_valid = PECross_237_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_238_multiply_io_input_io_actIn_bits_x_0 = PECross_237_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_238_multiply_io_input_io_actIn_bits_last = PECross_237_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_238_multiply_io_input_io_weiIn_valid = PECross_222_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_238_multiply_io_input_io_weiIn_bits_x_0 = PECross_222_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_238_multiply_io_input_io_weiIn_bits_last = PECross_222_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_238_multiply_io_input_io_actOut_ready = PECross_239_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_238_multiply_io_input_io_weiOut_ready = PECross_254_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_239_clock = clock;
  assign PECross_239_reset = rst;
  assign PECross_239_multiply_io_input_io_sumIn_valid = PECross_238_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_239_multiply_io_input_io_sumIn_bits_x_0 = PECross_238_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_239_multiply_io_input_io_sumIn_bits_last = PECross_238_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_239_multiply_io_input_io_sumOut_ready = io_sumOut_14_ready; // @[mac.scala 45:29]
  assign PECross_239_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_239_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_239_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_239_multiply_io_input_io_actIn_valid = PECross_238_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_239_multiply_io_input_io_actIn_bits_x_0 = PECross_238_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_239_multiply_io_input_io_actIn_bits_last = PECross_238_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_239_multiply_io_input_io_weiIn_valid = PECross_223_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_239_multiply_io_input_io_weiIn_bits_x_0 = PECross_223_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_239_multiply_io_input_io_weiIn_bits_last = PECross_223_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_239_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_239_multiply_io_input_io_weiOut_ready = PECross_255_multiply_io_input_io_weiIn_ready; // @[mac.scala 42:28]
  assign PECross_240_clock = clock;
  assign PECross_240_reset = rst;
  assign PECross_240_multiply_io_input_io_sumIn_valid = io_sumIn_15_valid; // @[mac.scala 33:28]
  assign PECross_240_multiply_io_input_io_sumIn_bits_x_0 = io_sumIn_15_bits_x_0; // @[mac.scala 33:28]
  assign PECross_240_multiply_io_input_io_sumIn_bits_last = io_sumIn_15_bits_last; // @[mac.scala 33:28]
  assign PECross_240_multiply_io_input_io_sumOut_ready = PECross_241_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_240_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_240_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_240_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_240_multiply_io_input_io_actIn_valid = io_actIn_15_valid; // @[mac.scala 32:28]
  assign PECross_240_multiply_io_input_io_actIn_bits_x_0 = io_actIn_15_bits_x_0; // @[mac.scala 32:28]
  assign PECross_240_multiply_io_input_io_actIn_bits_last = io_actIn_15_bits_last; // @[mac.scala 32:28]
  assign PECross_240_multiply_io_input_io_weiIn_valid = PECross_224_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_240_multiply_io_input_io_weiIn_bits_x_0 = PECross_224_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_240_multiply_io_input_io_weiIn_bits_last = PECross_224_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_240_multiply_io_input_io_actOut_ready = PECross_241_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_240_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_241_clock = clock;
  assign PECross_241_reset = rst;
  assign PECross_241_multiply_io_input_io_sumIn_valid = PECross_240_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_241_multiply_io_input_io_sumIn_bits_x_0 = PECross_240_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_241_multiply_io_input_io_sumIn_bits_last = PECross_240_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_241_multiply_io_input_io_sumOut_ready = PECross_242_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_241_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_241_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_241_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_241_multiply_io_input_io_actIn_valid = PECross_240_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_241_multiply_io_input_io_actIn_bits_x_0 = PECross_240_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_241_multiply_io_input_io_actIn_bits_last = PECross_240_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_241_multiply_io_input_io_weiIn_valid = PECross_225_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_241_multiply_io_input_io_weiIn_bits_x_0 = PECross_225_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_241_multiply_io_input_io_weiIn_bits_last = PECross_225_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_241_multiply_io_input_io_actOut_ready = PECross_242_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_241_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_242_clock = clock;
  assign PECross_242_reset = rst;
  assign PECross_242_multiply_io_input_io_sumIn_valid = PECross_241_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_242_multiply_io_input_io_sumIn_bits_x_0 = PECross_241_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_242_multiply_io_input_io_sumIn_bits_last = PECross_241_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_242_multiply_io_input_io_sumOut_ready = PECross_243_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_242_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_242_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_242_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_242_multiply_io_input_io_actIn_valid = PECross_241_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_242_multiply_io_input_io_actIn_bits_x_0 = PECross_241_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_242_multiply_io_input_io_actIn_bits_last = PECross_241_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_242_multiply_io_input_io_weiIn_valid = PECross_226_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_242_multiply_io_input_io_weiIn_bits_x_0 = PECross_226_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_242_multiply_io_input_io_weiIn_bits_last = PECross_226_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_242_multiply_io_input_io_actOut_ready = PECross_243_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_242_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_243_clock = clock;
  assign PECross_243_reset = rst;
  assign PECross_243_multiply_io_input_io_sumIn_valid = PECross_242_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_243_multiply_io_input_io_sumIn_bits_x_0 = PECross_242_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_243_multiply_io_input_io_sumIn_bits_last = PECross_242_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_243_multiply_io_input_io_sumOut_ready = PECross_244_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_243_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_243_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_243_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_243_multiply_io_input_io_actIn_valid = PECross_242_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_243_multiply_io_input_io_actIn_bits_x_0 = PECross_242_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_243_multiply_io_input_io_actIn_bits_last = PECross_242_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_243_multiply_io_input_io_weiIn_valid = PECross_227_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_243_multiply_io_input_io_weiIn_bits_x_0 = PECross_227_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_243_multiply_io_input_io_weiIn_bits_last = PECross_227_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_243_multiply_io_input_io_actOut_ready = PECross_244_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_243_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_244_clock = clock;
  assign PECross_244_reset = rst;
  assign PECross_244_multiply_io_input_io_sumIn_valid = PECross_243_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_244_multiply_io_input_io_sumIn_bits_x_0 = PECross_243_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_244_multiply_io_input_io_sumIn_bits_last = PECross_243_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_244_multiply_io_input_io_sumOut_ready = PECross_245_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_244_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_244_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_244_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_244_multiply_io_input_io_actIn_valid = PECross_243_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_244_multiply_io_input_io_actIn_bits_x_0 = PECross_243_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_244_multiply_io_input_io_actIn_bits_last = PECross_243_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_244_multiply_io_input_io_weiIn_valid = PECross_228_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_244_multiply_io_input_io_weiIn_bits_x_0 = PECross_228_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_244_multiply_io_input_io_weiIn_bits_last = PECross_228_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_244_multiply_io_input_io_actOut_ready = PECross_245_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_244_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_245_clock = clock;
  assign PECross_245_reset = rst;
  assign PECross_245_multiply_io_input_io_sumIn_valid = PECross_244_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_245_multiply_io_input_io_sumIn_bits_x_0 = PECross_244_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_245_multiply_io_input_io_sumIn_bits_last = PECross_244_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_245_multiply_io_input_io_sumOut_ready = PECross_246_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_245_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_245_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_245_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_245_multiply_io_input_io_actIn_valid = PECross_244_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_245_multiply_io_input_io_actIn_bits_x_0 = PECross_244_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_245_multiply_io_input_io_actIn_bits_last = PECross_244_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_245_multiply_io_input_io_weiIn_valid = PECross_229_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_245_multiply_io_input_io_weiIn_bits_x_0 = PECross_229_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_245_multiply_io_input_io_weiIn_bits_last = PECross_229_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_245_multiply_io_input_io_actOut_ready = PECross_246_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_245_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_246_clock = clock;
  assign PECross_246_reset = rst;
  assign PECross_246_multiply_io_input_io_sumIn_valid = PECross_245_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_246_multiply_io_input_io_sumIn_bits_x_0 = PECross_245_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_246_multiply_io_input_io_sumIn_bits_last = PECross_245_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_246_multiply_io_input_io_sumOut_ready = PECross_247_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_246_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_246_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_246_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_246_multiply_io_input_io_actIn_valid = PECross_245_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_246_multiply_io_input_io_actIn_bits_x_0 = PECross_245_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_246_multiply_io_input_io_actIn_bits_last = PECross_245_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_246_multiply_io_input_io_weiIn_valid = PECross_230_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_246_multiply_io_input_io_weiIn_bits_x_0 = PECross_230_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_246_multiply_io_input_io_weiIn_bits_last = PECross_230_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_246_multiply_io_input_io_actOut_ready = PECross_247_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_246_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_247_clock = clock;
  assign PECross_247_reset = rst;
  assign PECross_247_multiply_io_input_io_sumIn_valid = PECross_246_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_247_multiply_io_input_io_sumIn_bits_x_0 = PECross_246_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_247_multiply_io_input_io_sumIn_bits_last = PECross_246_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_247_multiply_io_input_io_sumOut_ready = PECross_248_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_247_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_247_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_247_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_247_multiply_io_input_io_actIn_valid = PECross_246_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_247_multiply_io_input_io_actIn_bits_x_0 = PECross_246_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_247_multiply_io_input_io_actIn_bits_last = PECross_246_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_247_multiply_io_input_io_weiIn_valid = PECross_231_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_247_multiply_io_input_io_weiIn_bits_x_0 = PECross_231_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_247_multiply_io_input_io_weiIn_bits_last = PECross_231_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_247_multiply_io_input_io_actOut_ready = PECross_248_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_247_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_248_clock = clock;
  assign PECross_248_reset = rst;
  assign PECross_248_multiply_io_input_io_sumIn_valid = PECross_247_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_248_multiply_io_input_io_sumIn_bits_x_0 = PECross_247_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_248_multiply_io_input_io_sumIn_bits_last = PECross_247_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_248_multiply_io_input_io_sumOut_ready = PECross_249_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_248_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_248_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_248_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_248_multiply_io_input_io_actIn_valid = PECross_247_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_248_multiply_io_input_io_actIn_bits_x_0 = PECross_247_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_248_multiply_io_input_io_actIn_bits_last = PECross_247_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_248_multiply_io_input_io_weiIn_valid = PECross_232_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_248_multiply_io_input_io_weiIn_bits_x_0 = PECross_232_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_248_multiply_io_input_io_weiIn_bits_last = PECross_232_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_248_multiply_io_input_io_actOut_ready = PECross_249_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_248_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_249_clock = clock;
  assign PECross_249_reset = rst;
  assign PECross_249_multiply_io_input_io_sumIn_valid = PECross_248_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_249_multiply_io_input_io_sumIn_bits_x_0 = PECross_248_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_249_multiply_io_input_io_sumIn_bits_last = PECross_248_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_249_multiply_io_input_io_sumOut_ready = PECross_250_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_249_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_249_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_249_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_249_multiply_io_input_io_actIn_valid = PECross_248_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_249_multiply_io_input_io_actIn_bits_x_0 = PECross_248_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_249_multiply_io_input_io_actIn_bits_last = PECross_248_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_249_multiply_io_input_io_weiIn_valid = PECross_233_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_249_multiply_io_input_io_weiIn_bits_x_0 = PECross_233_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_249_multiply_io_input_io_weiIn_bits_last = PECross_233_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_249_multiply_io_input_io_actOut_ready = PECross_250_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_249_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_250_clock = clock;
  assign PECross_250_reset = rst;
  assign PECross_250_multiply_io_input_io_sumIn_valid = PECross_249_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_250_multiply_io_input_io_sumIn_bits_x_0 = PECross_249_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_250_multiply_io_input_io_sumIn_bits_last = PECross_249_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_250_multiply_io_input_io_sumOut_ready = PECross_251_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_250_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_250_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_250_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_250_multiply_io_input_io_actIn_valid = PECross_249_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_250_multiply_io_input_io_actIn_bits_x_0 = PECross_249_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_250_multiply_io_input_io_actIn_bits_last = PECross_249_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_250_multiply_io_input_io_weiIn_valid = PECross_234_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_250_multiply_io_input_io_weiIn_bits_x_0 = PECross_234_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_250_multiply_io_input_io_weiIn_bits_last = PECross_234_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_250_multiply_io_input_io_actOut_ready = PECross_251_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_250_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_251_clock = clock;
  assign PECross_251_reset = rst;
  assign PECross_251_multiply_io_input_io_sumIn_valid = PECross_250_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_251_multiply_io_input_io_sumIn_bits_x_0 = PECross_250_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_251_multiply_io_input_io_sumIn_bits_last = PECross_250_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_251_multiply_io_input_io_sumOut_ready = PECross_252_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_251_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_251_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_251_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_251_multiply_io_input_io_actIn_valid = PECross_250_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_251_multiply_io_input_io_actIn_bits_x_0 = PECross_250_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_251_multiply_io_input_io_actIn_bits_last = PECross_250_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_251_multiply_io_input_io_weiIn_valid = PECross_235_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_251_multiply_io_input_io_weiIn_bits_x_0 = PECross_235_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_251_multiply_io_input_io_weiIn_bits_last = PECross_235_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_251_multiply_io_input_io_actOut_ready = PECross_252_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_251_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_252_clock = clock;
  assign PECross_252_reset = rst;
  assign PECross_252_multiply_io_input_io_sumIn_valid = PECross_251_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_252_multiply_io_input_io_sumIn_bits_x_0 = PECross_251_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_252_multiply_io_input_io_sumIn_bits_last = PECross_251_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_252_multiply_io_input_io_sumOut_ready = PECross_253_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_252_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_252_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_252_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_252_multiply_io_input_io_actIn_valid = PECross_251_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_252_multiply_io_input_io_actIn_bits_x_0 = PECross_251_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_252_multiply_io_input_io_actIn_bits_last = PECross_251_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_252_multiply_io_input_io_weiIn_valid = PECross_236_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_252_multiply_io_input_io_weiIn_bits_x_0 = PECross_236_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_252_multiply_io_input_io_weiIn_bits_last = PECross_236_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_252_multiply_io_input_io_actOut_ready = PECross_253_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_252_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_253_clock = clock;
  assign PECross_253_reset = rst;
  assign PECross_253_multiply_io_input_io_sumIn_valid = PECross_252_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_253_multiply_io_input_io_sumIn_bits_x_0 = PECross_252_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_253_multiply_io_input_io_sumIn_bits_last = PECross_252_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_253_multiply_io_input_io_sumOut_ready = PECross_254_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_253_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_253_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_253_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_253_multiply_io_input_io_actIn_valid = PECross_252_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_253_multiply_io_input_io_actIn_bits_x_0 = PECross_252_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_253_multiply_io_input_io_actIn_bits_last = PECross_252_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_253_multiply_io_input_io_weiIn_valid = PECross_237_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_253_multiply_io_input_io_weiIn_bits_x_0 = PECross_237_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_253_multiply_io_input_io_weiIn_bits_last = PECross_237_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_253_multiply_io_input_io_actOut_ready = PECross_254_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_253_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_254_clock = clock;
  assign PECross_254_reset = rst;
  assign PECross_254_multiply_io_input_io_sumIn_valid = PECross_253_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_254_multiply_io_input_io_sumIn_bits_x_0 = PECross_253_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_254_multiply_io_input_io_sumIn_bits_last = PECross_253_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_254_multiply_io_input_io_sumOut_ready = PECross_255_multiply_io_input_io_sumIn_ready; // @[mac.scala 37:28]
  assign PECross_254_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_254_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_254_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_254_multiply_io_input_io_actIn_valid = PECross_253_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_254_multiply_io_input_io_actIn_bits_x_0 = PECross_253_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_254_multiply_io_input_io_actIn_bits_last = PECross_253_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_254_multiply_io_input_io_weiIn_valid = PECross_238_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_254_multiply_io_input_io_weiIn_bits_x_0 = PECross_238_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_254_multiply_io_input_io_weiIn_bits_last = PECross_238_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_254_multiply_io_input_io_actOut_ready = PECross_255_multiply_io_input_io_actIn_ready; // @[mac.scala 36:28]
  assign PECross_254_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
  assign PECross_255_clock = clock;
  assign PECross_255_reset = rst;
  assign PECross_255_multiply_io_input_io_sumIn_valid = PECross_254_multiply_io_input_io_sumOut_valid; // @[mac.scala 37:28]
  assign PECross_255_multiply_io_input_io_sumIn_bits_x_0 = PECross_254_multiply_io_input_io_sumOut_bits_x_0; // @[mac.scala 37:28]
  assign PECross_255_multiply_io_input_io_sumIn_bits_last = PECross_254_multiply_io_input_io_sumOut_bits_last; // @[mac.scala 37:28]
  assign PECross_255_multiply_io_input_io_sumOut_ready = io_sumOut_15_ready; // @[mac.scala 45:29]
  assign PECross_255_multiply_io_input_io_statSel = io_statSel; // @[mac.scala 53:26]
  assign PECross_255_multiply_io_input_io_weiEn = io_weiEn; // @[mac.scala 55:24]
  assign PECross_255_multiply_io_input_io_actEn = io_actEn; // @[mac.scala 54:24]
  assign PECross_255_multiply_io_input_io_actIn_valid = PECross_254_multiply_io_input_io_actOut_valid; // @[mac.scala 36:28]
  assign PECross_255_multiply_io_input_io_actIn_bits_x_0 = PECross_254_multiply_io_input_io_actOut_bits_x_0; // @[mac.scala 36:28]
  assign PECross_255_multiply_io_input_io_actIn_bits_last = PECross_254_multiply_io_input_io_actOut_bits_last; // @[mac.scala 36:28]
  assign PECross_255_multiply_io_input_io_weiIn_valid = PECross_239_multiply_io_input_io_weiOut_valid; // @[mac.scala 42:28]
  assign PECross_255_multiply_io_input_io_weiIn_bits_x_0 = PECross_239_multiply_io_input_io_weiOut_bits_x_0; // @[mac.scala 42:28]
  assign PECross_255_multiply_io_input_io_weiIn_bits_last = PECross_239_multiply_io_input_io_weiOut_bits_last; // @[mac.scala 42:28]
  assign PECross_255_multiply_io_input_io_actOut_ready = io_actOutReady; // @[mac.scala 44:35]
  assign PECross_255_multiply_io_input_io_weiOut_ready = io_weiOutReady; // @[mac.scala 48:35]
endmodule
